`timescale  1ns/1ns
 
module tb_result4_2x2;
 
parameter  T = 2; // 时钟周期 ns
 
reg          clk; //input 
reg          rst_n; //input 
reg  [7:0]  dq_i; //input 
reg  [10:0]  xpos; //input 
reg  [10:0]  ypos; //input 
wire [4:0]  digit; //output 

// *******************************************************************************
// ** main
// *******************************************************************************

initial begin
   clk      =1'b0;
   rst_n      =1'b0;
 
   #T //1 start
// 20.0 ns
   rst_n      =1'b1;
 
   #T//
   xpos = 211;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 214;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 215;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 216;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 217;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 218;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 219;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 220;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 221;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 222;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 223;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 224;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 225;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 226;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 227;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 228;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 229;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 230;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 231;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 232;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 233;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 234;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 235;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 236;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 237;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 238;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 239;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 240;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 241;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 242;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 243;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 244;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 245;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 246;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 247;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 248;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 249;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 250;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 251;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 252;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 253;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 254;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 255;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 256;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 257;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 258;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 259;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 260;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 261;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 262;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 263;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 264;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 265;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 266;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 267;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 268;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 269;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 107;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 214;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 215;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 216;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 217;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 218;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 219;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 220;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 221;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 222;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 223;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 224;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 225;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 226;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 227;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 228;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 229;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 230;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 231;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 232;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 233;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 234;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 235;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 236;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 237;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 238;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 239;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 240;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 241;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 242;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 243;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 244;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 245;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 246;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 247;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 248;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 249;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 250;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 251;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 252;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 253;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 254;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 255;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 256;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 257;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 258;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 259;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 260;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 261;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 262;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 263;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 264;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 265;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 266;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 267;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 268;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 269;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 108;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 109;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 109;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 109;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 109;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 109;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 110;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 110;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 110;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 110;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 110;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 111;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 111;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 111;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 111;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 111;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 112;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 112;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 112;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 112;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 112;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 113;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 113;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 113;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 113;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 113;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 114;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 114;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 114;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 114;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 114;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 115;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 115;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 115;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 115;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 115;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 116;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 116;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 116;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 116;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 116;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 117;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 117;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 117;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 117;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 117;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 118;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 118;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 118;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 118;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 118;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 119;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 119;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 119;
   dq_i = 50;
 
   #T//
   xpos = 234;
   ypos = 119;
   dq_i = 50;
 
   #T//
   xpos = 235;
   ypos = 119;
   dq_i = 224;
 
   #T//
   xpos = 236;
   ypos = 119;
   dq_i = 224;
 
   #T//
   xpos = 237;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 119;
   dq_i = 70;
 
   #T//
   xpos = 252;
   ypos = 119;
   dq_i = 70;
 
   #T//
   xpos = 253;
   ypos = 119;
   dq_i = 29;
 
   #T//
   xpos = 254;
   ypos = 119;
   dq_i = 29;
 
   #T//
   xpos = 255;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 119;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 119;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 119;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 120;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 120;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 120;
   dq_i = 50;
 
   #T//
   xpos = 234;
   ypos = 120;
   dq_i = 50;
 
   #T//
   xpos = 235;
   ypos = 120;
   dq_i = 224;
 
   #T//
   xpos = 236;
   ypos = 120;
   dq_i = 224;
 
   #T//
   xpos = 237;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 120;
   dq_i = 70;
 
   #T//
   xpos = 252;
   ypos = 120;
   dq_i = 70;
 
   #T//
   xpos = 253;
   ypos = 120;
   dq_i = 29;
 
   #T//
   xpos = 254;
   ypos = 120;
   dq_i = 29;
 
   #T//
   xpos = 255;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 120;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 120;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 120;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 121;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 121;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 121;
   dq_i = 121;
 
   #T//
   xpos = 234;
   ypos = 121;
   dq_i = 121;
 
   #T//
   xpos = 235;
   ypos = 121;
   dq_i = 231;
 
   #T//
   xpos = 236;
   ypos = 121;
   dq_i = 231;
 
   #T//
   xpos = 237;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 121;
   dq_i = 148;
 
   #T//
   xpos = 252;
   ypos = 121;
   dq_i = 148;
 
   #T//
   xpos = 253;
   ypos = 121;
   dq_i = 168;
 
   #T//
   xpos = 254;
   ypos = 121;
   dq_i = 168;
 
   #T//
   xpos = 255;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 121;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 121;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 121;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 122;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 122;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 122;
   dq_i = 121;
 
   #T//
   xpos = 234;
   ypos = 122;
   dq_i = 121;
 
   #T//
   xpos = 235;
   ypos = 122;
   dq_i = 231;
 
   #T//
   xpos = 236;
   ypos = 122;
   dq_i = 231;
 
   #T//
   xpos = 237;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 122;
   dq_i = 148;
 
   #T//
   xpos = 252;
   ypos = 122;
   dq_i = 148;
 
   #T//
   xpos = 253;
   ypos = 122;
   dq_i = 168;
 
   #T//
   xpos = 254;
   ypos = 122;
   dq_i = 168;
 
   #T//
   xpos = 255;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 122;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 122;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 122;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 123;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 123;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 123;
   dq_i = 4;
 
   #T//
   xpos = 232;
   ypos = 123;
   dq_i = 4;
 
   #T//
   xpos = 233;
   ypos = 123;
   dq_i = 195;
 
   #T//
   xpos = 234;
   ypos = 123;
   dq_i = 195;
 
   #T//
   xpos = 235;
   ypos = 123;
   dq_i = 231;
 
   #T//
   xpos = 236;
   ypos = 123;
   dq_i = 231;
 
   #T//
   xpos = 237;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 123;
   dq_i = 96;
 
   #T//
   xpos = 252;
   ypos = 123;
   dq_i = 96;
 
   #T//
   xpos = 253;
   ypos = 123;
   dq_i = 210;
 
   #T//
   xpos = 254;
   ypos = 123;
   dq_i = 210;
 
   #T//
   xpos = 255;
   ypos = 123;
   dq_i = 11;
 
   #T//
   xpos = 256;
   ypos = 123;
   dq_i = 11;
 
   #T//
   xpos = 257;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 123;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 123;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 123;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 124;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 124;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 124;
   dq_i = 4;
 
   #T//
   xpos = 232;
   ypos = 124;
   dq_i = 4;
 
   #T//
   xpos = 233;
   ypos = 124;
   dq_i = 195;
 
   #T//
   xpos = 234;
   ypos = 124;
   dq_i = 195;
 
   #T//
   xpos = 235;
   ypos = 124;
   dq_i = 231;
 
   #T//
   xpos = 236;
   ypos = 124;
   dq_i = 231;
 
   #T//
   xpos = 237;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 124;
   dq_i = 96;
 
   #T//
   xpos = 252;
   ypos = 124;
   dq_i = 96;
 
   #T//
   xpos = 253;
   ypos = 124;
   dq_i = 210;
 
   #T//
   xpos = 254;
   ypos = 124;
   dq_i = 210;
 
   #T//
   xpos = 255;
   ypos = 124;
   dq_i = 11;
 
   #T//
   xpos = 256;
   ypos = 124;
   dq_i = 11;
 
   #T//
   xpos = 257;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 124;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 124;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 124;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 125;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 125;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 125;
   dq_i = 69;
 
   #T//
   xpos = 232;
   ypos = 125;
   dq_i = 69;
 
   #T//
   xpos = 233;
   ypos = 125;
   dq_i = 252;
 
   #T//
   xpos = 234;
   ypos = 125;
   dq_i = 252;
 
   #T//
   xpos = 235;
   ypos = 125;
   dq_i = 134;
 
   #T//
   xpos = 236;
   ypos = 125;
   dq_i = 134;
 
   #T//
   xpos = 237;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 125;
   dq_i = 114;
 
   #T//
   xpos = 252;
   ypos = 125;
   dq_i = 114;
 
   #T//
   xpos = 253;
   ypos = 125;
   dq_i = 252;
 
   #T//
   xpos = 254;
   ypos = 125;
   dq_i = 252;
 
   #T//
   xpos = 255;
   ypos = 125;
   dq_i = 21;
 
   #T//
   xpos = 256;
   ypos = 125;
   dq_i = 21;
 
   #T//
   xpos = 257;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 125;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 125;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 125;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 126;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 126;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 126;
   dq_i = 69;
 
   #T//
   xpos = 232;
   ypos = 126;
   dq_i = 69;
 
   #T//
   xpos = 233;
   ypos = 126;
   dq_i = 252;
 
   #T//
   xpos = 234;
   ypos = 126;
   dq_i = 252;
 
   #T//
   xpos = 235;
   ypos = 126;
   dq_i = 134;
 
   #T//
   xpos = 236;
   ypos = 126;
   dq_i = 134;
 
   #T//
   xpos = 237;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 126;
   dq_i = 114;
 
   #T//
   xpos = 252;
   ypos = 126;
   dq_i = 114;
 
   #T//
   xpos = 253;
   ypos = 126;
   dq_i = 252;
 
   #T//
   xpos = 254;
   ypos = 126;
   dq_i = 252;
 
   #T//
   xpos = 255;
   ypos = 126;
   dq_i = 21;
 
   #T//
   xpos = 256;
   ypos = 126;
   dq_i = 21;
 
   #T//
   xpos = 257;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 126;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 126;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 126;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 127;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 127;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 127;
   dq_i = 45;
 
   #T//
   xpos = 230;
   ypos = 127;
   dq_i = 45;
 
   #T//
   xpos = 231;
   ypos = 127;
   dq_i = 236;
 
   #T//
   xpos = 232;
   ypos = 127;
   dq_i = 236;
 
   #T//
   xpos = 233;
   ypos = 127;
   dq_i = 217;
 
   #T//
   xpos = 234;
   ypos = 127;
   dq_i = 217;
 
   #T//
   xpos = 235;
   ypos = 127;
   dq_i = 12;
 
   #T//
   xpos = 236;
   ypos = 127;
   dq_i = 12;
 
   #T//
   xpos = 237;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 127;
   dq_i = 192;
 
   #T//
   xpos = 252;
   ypos = 127;
   dq_i = 192;
 
   #T//
   xpos = 253;
   ypos = 127;
   dq_i = 252;
 
   #T//
   xpos = 254;
   ypos = 127;
   dq_i = 252;
 
   #T//
   xpos = 255;
   ypos = 127;
   dq_i = 21;
 
   #T//
   xpos = 256;
   ypos = 127;
   dq_i = 21;
 
   #T//
   xpos = 257;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 127;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 127;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 127;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 128;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 128;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 128;
   dq_i = 45;
 
   #T//
   xpos = 230;
   ypos = 128;
   dq_i = 45;
 
   #T//
   xpos = 231;
   ypos = 128;
   dq_i = 236;
 
   #T//
   xpos = 232;
   ypos = 128;
   dq_i = 236;
 
   #T//
   xpos = 233;
   ypos = 128;
   dq_i = 217;
 
   #T//
   xpos = 234;
   ypos = 128;
   dq_i = 217;
 
   #T//
   xpos = 235;
   ypos = 128;
   dq_i = 12;
 
   #T//
   xpos = 236;
   ypos = 128;
   dq_i = 12;
 
   #T//
   xpos = 237;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 128;
   dq_i = 192;
 
   #T//
   xpos = 252;
   ypos = 128;
   dq_i = 192;
 
   #T//
   xpos = 253;
   ypos = 128;
   dq_i = 252;
 
   #T//
   xpos = 254;
   ypos = 128;
   dq_i = 252;
 
   #T//
   xpos = 255;
   ypos = 128;
   dq_i = 21;
 
   #T//
   xpos = 256;
   ypos = 128;
   dq_i = 21;
 
   #T//
   xpos = 257;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 128;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 128;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 128;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 129;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 129;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 129;
   dq_i = 168;
 
   #T//
   xpos = 230;
   ypos = 129;
   dq_i = 168;
 
   #T//
   xpos = 231;
   ypos = 129;
   dq_i = 247;
 
   #T//
   xpos = 232;
   ypos = 129;
   dq_i = 247;
 
   #T//
   xpos = 233;
   ypos = 129;
   dq_i = 53;
 
   #T//
   xpos = 234;
   ypos = 129;
   dq_i = 53;
 
   #T//
   xpos = 235;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 129;
   dq_i = 18;
 
   #T//
   xpos = 250;
   ypos = 129;
   dq_i = 18;
 
   #T//
   xpos = 251;
   ypos = 129;
   dq_i = 255;
 
   #T//
   xpos = 252;
   ypos = 129;
   dq_i = 255;
 
   #T//
   xpos = 253;
   ypos = 129;
   dq_i = 253;
 
   #T//
   xpos = 254;
   ypos = 129;
   dq_i = 253;
 
   #T//
   xpos = 255;
   ypos = 129;
   dq_i = 21;
 
   #T//
   xpos = 256;
   ypos = 129;
   dq_i = 21;
 
   #T//
   xpos = 257;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 129;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 129;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 129;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 130;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 130;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 130;
   dq_i = 168;
 
   #T//
   xpos = 230;
   ypos = 130;
   dq_i = 168;
 
   #T//
   xpos = 231;
   ypos = 130;
   dq_i = 247;
 
   #T//
   xpos = 232;
   ypos = 130;
   dq_i = 247;
 
   #T//
   xpos = 233;
   ypos = 130;
   dq_i = 53;
 
   #T//
   xpos = 234;
   ypos = 130;
   dq_i = 53;
 
   #T//
   xpos = 235;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 130;
   dq_i = 18;
 
   #T//
   xpos = 250;
   ypos = 130;
   dq_i = 18;
 
   #T//
   xpos = 251;
   ypos = 130;
   dq_i = 255;
 
   #T//
   xpos = 252;
   ypos = 130;
   dq_i = 255;
 
   #T//
   xpos = 253;
   ypos = 130;
   dq_i = 253;
 
   #T//
   xpos = 254;
   ypos = 130;
   dq_i = 253;
 
   #T//
   xpos = 255;
   ypos = 130;
   dq_i = 21;
 
   #T//
   xpos = 256;
   ypos = 130;
   dq_i = 21;
 
   #T//
   xpos = 257;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 130;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 130;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 130;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 131;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 131;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 131;
   dq_i = 84;
 
   #T//
   xpos = 228;
   ypos = 131;
   dq_i = 84;
 
   #T//
   xpos = 229;
   ypos = 131;
   dq_i = 242;
 
   #T//
   xpos = 230;
   ypos = 131;
   dq_i = 242;
 
   #T//
   xpos = 231;
   ypos = 131;
   dq_i = 211;
 
   #T//
   xpos = 232;
   ypos = 131;
   dq_i = 211;
 
   #T//
   xpos = 233;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 131;
   dq_i = 141;
 
   #T//
   xpos = 250;
   ypos = 131;
   dq_i = 141;
 
   #T//
   xpos = 251;
   ypos = 131;
   dq_i = 253;
 
   #T//
   xpos = 252;
   ypos = 131;
   dq_i = 253;
 
   #T//
   xpos = 253;
   ypos = 131;
   dq_i = 189;
 
   #T//
   xpos = 254;
   ypos = 131;
   dq_i = 189;
 
   #T//
   xpos = 255;
   ypos = 131;
   dq_i = 5;
 
   #T//
   xpos = 256;
   ypos = 131;
   dq_i = 5;
 
   #T//
   xpos = 257;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 131;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 131;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 131;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 132;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 132;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 132;
   dq_i = 84;
 
   #T//
   xpos = 228;
   ypos = 132;
   dq_i = 84;
 
   #T//
   xpos = 229;
   ypos = 132;
   dq_i = 242;
 
   #T//
   xpos = 230;
   ypos = 132;
   dq_i = 242;
 
   #T//
   xpos = 231;
   ypos = 132;
   dq_i = 211;
 
   #T//
   xpos = 232;
   ypos = 132;
   dq_i = 211;
 
   #T//
   xpos = 233;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 132;
   dq_i = 141;
 
   #T//
   xpos = 250;
   ypos = 132;
   dq_i = 141;
 
   #T//
   xpos = 251;
   ypos = 132;
   dq_i = 253;
 
   #T//
   xpos = 252;
   ypos = 132;
   dq_i = 253;
 
   #T//
   xpos = 253;
   ypos = 132;
   dq_i = 189;
 
   #T//
   xpos = 254;
   ypos = 132;
   dq_i = 189;
 
   #T//
   xpos = 255;
   ypos = 132;
   dq_i = 5;
 
   #T//
   xpos = 256;
   ypos = 132;
   dq_i = 5;
 
   #T//
   xpos = 257;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 132;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 132;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 132;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 133;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 133;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 133;
   dq_i = 169;
 
   #T//
   xpos = 228;
   ypos = 133;
   dq_i = 169;
 
   #T//
   xpos = 229;
   ypos = 133;
   dq_i = 252;
 
   #T//
   xpos = 230;
   ypos = 133;
   dq_i = 252;
 
   #T//
   xpos = 231;
   ypos = 133;
   dq_i = 106;
 
   #T//
   xpos = 232;
   ypos = 133;
   dq_i = 106;
 
   #T//
   xpos = 233;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 133;
   dq_i = 32;
 
   #T//
   xpos = 248;
   ypos = 133;
   dq_i = 32;
 
   #T//
   xpos = 249;
   ypos = 133;
   dq_i = 232;
 
   #T//
   xpos = 250;
   ypos = 133;
   dq_i = 232;
 
   #T//
   xpos = 251;
   ypos = 133;
   dq_i = 250;
 
   #T//
   xpos = 252;
   ypos = 133;
   dq_i = 250;
 
   #T//
   xpos = 253;
   ypos = 133;
   dq_i = 66;
 
   #T//
   xpos = 254;
   ypos = 133;
   dq_i = 66;
 
   #T//
   xpos = 255;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 133;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 133;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 133;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 134;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 134;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 134;
   dq_i = 169;
 
   #T//
   xpos = 228;
   ypos = 134;
   dq_i = 169;
 
   #T//
   xpos = 229;
   ypos = 134;
   dq_i = 252;
 
   #T//
   xpos = 230;
   ypos = 134;
   dq_i = 252;
 
   #T//
   xpos = 231;
   ypos = 134;
   dq_i = 106;
 
   #T//
   xpos = 232;
   ypos = 134;
   dq_i = 106;
 
   #T//
   xpos = 233;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 134;
   dq_i = 32;
 
   #T//
   xpos = 248;
   ypos = 134;
   dq_i = 32;
 
   #T//
   xpos = 249;
   ypos = 134;
   dq_i = 232;
 
   #T//
   xpos = 250;
   ypos = 134;
   dq_i = 232;
 
   #T//
   xpos = 251;
   ypos = 134;
   dq_i = 250;
 
   #T//
   xpos = 252;
   ypos = 134;
   dq_i = 250;
 
   #T//
   xpos = 253;
   ypos = 134;
   dq_i = 66;
 
   #T//
   xpos = 254;
   ypos = 134;
   dq_i = 66;
 
   #T//
   xpos = 255;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 134;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 134;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 134;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 135;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 135;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 135;
   dq_i = 15;
 
   #T//
   xpos = 226;
   ypos = 135;
   dq_i = 15;
 
   #T//
   xpos = 227;
   ypos = 135;
   dq_i = 225;
 
   #T//
   xpos = 228;
   ypos = 135;
   dq_i = 225;
 
   #T//
   xpos = 229;
   ypos = 135;
   dq_i = 252;
 
   #T//
   xpos = 230;
   ypos = 135;
   dq_i = 252;
 
   #T//
   xpos = 231;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 135;
   dq_i = 134;
 
   #T//
   xpos = 248;
   ypos = 135;
   dq_i = 134;
 
   #T//
   xpos = 249;
   ypos = 135;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 135;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 135;
   dq_i = 211;
 
   #T//
   xpos = 252;
   ypos = 135;
   dq_i = 211;
 
   #T//
   xpos = 253;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 135;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 135;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 135;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 136;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 136;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 136;
   dq_i = 15;
 
   #T//
   xpos = 226;
   ypos = 136;
   dq_i = 15;
 
   #T//
   xpos = 227;
   ypos = 136;
   dq_i = 225;
 
   #T//
   xpos = 228;
   ypos = 136;
   dq_i = 225;
 
   #T//
   xpos = 229;
   ypos = 136;
   dq_i = 252;
 
   #T//
   xpos = 230;
   ypos = 136;
   dq_i = 252;
 
   #T//
   xpos = 231;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 136;
   dq_i = 134;
 
   #T//
   xpos = 248;
   ypos = 136;
   dq_i = 134;
 
   #T//
   xpos = 249;
   ypos = 136;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 136;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 136;
   dq_i = 211;
 
   #T//
   xpos = 252;
   ypos = 136;
   dq_i = 211;
 
   #T//
   xpos = 253;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 136;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 136;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 136;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 137;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 137;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 137;
   dq_i = 22;
 
   #T//
   xpos = 226;
   ypos = 137;
   dq_i = 22;
 
   #T//
   xpos = 227;
   ypos = 137;
   dq_i = 252;
 
   #T//
   xpos = 228;
   ypos = 137;
   dq_i = 252;
 
   #T//
   xpos = 229;
   ypos = 137;
   dq_i = 164;
 
   #T//
   xpos = 230;
   ypos = 137;
   dq_i = 164;
 
   #T//
   xpos = 231;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 137;
   dq_i = 169;
 
   #T//
   xpos = 248;
   ypos = 137;
   dq_i = 169;
 
   #T//
   xpos = 249;
   ypos = 137;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 137;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 137;
   dq_i = 167;
 
   #T//
   xpos = 252;
   ypos = 137;
   dq_i = 167;
 
   #T//
   xpos = 253;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 137;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 137;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 137;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 138;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 138;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 138;
   dq_i = 22;
 
   #T//
   xpos = 226;
   ypos = 138;
   dq_i = 22;
 
   #T//
   xpos = 227;
   ypos = 138;
   dq_i = 252;
 
   #T//
   xpos = 228;
   ypos = 138;
   dq_i = 252;
 
   #T//
   xpos = 229;
   ypos = 138;
   dq_i = 164;
 
   #T//
   xpos = 230;
   ypos = 138;
   dq_i = 164;
 
   #T//
   xpos = 231;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 138;
   dq_i = 169;
 
   #T//
   xpos = 248;
   ypos = 138;
   dq_i = 169;
 
   #T//
   xpos = 249;
   ypos = 138;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 138;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 138;
   dq_i = 167;
 
   #T//
   xpos = 252;
   ypos = 138;
   dq_i = 167;
 
   #T//
   xpos = 253;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 138;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 138;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 138;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 139;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 139;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 139;
   dq_i = 9;
 
   #T//
   xpos = 226;
   ypos = 139;
   dq_i = 9;
 
   #T//
   xpos = 227;
   ypos = 139;
   dq_i = 204;
 
   #T//
   xpos = 228;
   ypos = 139;
   dq_i = 204;
 
   #T//
   xpos = 229;
   ypos = 139;
   dq_i = 209;
 
   #T//
   xpos = 230;
   ypos = 139;
   dq_i = 209;
 
   #T//
   xpos = 231;
   ypos = 139;
   dq_i = 18;
 
   #T//
   xpos = 232;
   ypos = 139;
   dq_i = 18;
 
   #T//
   xpos = 233;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 139;
   dq_i = 22;
 
   #T//
   xpos = 246;
   ypos = 139;
   dq_i = 22;
 
   #T//
   xpos = 247;
   ypos = 139;
   dq_i = 253;
 
   #T//
   xpos = 248;
   ypos = 139;
   dq_i = 253;
 
   #T//
   xpos = 249;
   ypos = 139;
   dq_i = 253;
 
   #T//
   xpos = 250;
   ypos = 139;
   dq_i = 253;
 
   #T//
   xpos = 251;
   ypos = 139;
   dq_i = 107;
 
   #T//
   xpos = 252;
   ypos = 139;
   dq_i = 107;
 
   #T//
   xpos = 253;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 139;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 139;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 139;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 140;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 140;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 140;
   dq_i = 9;
 
   #T//
   xpos = 226;
   ypos = 140;
   dq_i = 9;
 
   #T//
   xpos = 227;
   ypos = 140;
   dq_i = 204;
 
   #T//
   xpos = 228;
   ypos = 140;
   dq_i = 204;
 
   #T//
   xpos = 229;
   ypos = 140;
   dq_i = 209;
 
   #T//
   xpos = 230;
   ypos = 140;
   dq_i = 209;
 
   #T//
   xpos = 231;
   ypos = 140;
   dq_i = 18;
 
   #T//
   xpos = 232;
   ypos = 140;
   dq_i = 18;
 
   #T//
   xpos = 233;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 140;
   dq_i = 22;
 
   #T//
   xpos = 246;
   ypos = 140;
   dq_i = 22;
 
   #T//
   xpos = 247;
   ypos = 140;
   dq_i = 253;
 
   #T//
   xpos = 248;
   ypos = 140;
   dq_i = 253;
 
   #T//
   xpos = 249;
   ypos = 140;
   dq_i = 253;
 
   #T//
   xpos = 250;
   ypos = 140;
   dq_i = 253;
 
   #T//
   xpos = 251;
   ypos = 140;
   dq_i = 107;
 
   #T//
   xpos = 252;
   ypos = 140;
   dq_i = 107;
 
   #T//
   xpos = 253;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 140;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 140;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 140;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 141;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 141;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 141;
   dq_i = 169;
 
   #T//
   xpos = 228;
   ypos = 141;
   dq_i = 169;
 
   #T//
   xpos = 229;
   ypos = 141;
   dq_i = 252;
 
   #T//
   xpos = 230;
   ypos = 141;
   dq_i = 252;
 
   #T//
   xpos = 231;
   ypos = 141;
   dq_i = 199;
 
   #T//
   xpos = 232;
   ypos = 141;
   dq_i = 199;
 
   #T//
   xpos = 233;
   ypos = 141;
   dq_i = 85;
 
   #T//
   xpos = 234;
   ypos = 141;
   dq_i = 85;
 
   #T//
   xpos = 235;
   ypos = 141;
   dq_i = 85;
 
   #T//
   xpos = 236;
   ypos = 141;
   dq_i = 85;
 
   #T//
   xpos = 237;
   ypos = 141;
   dq_i = 85;
 
   #T//
   xpos = 238;
   ypos = 141;
   dq_i = 85;
 
   #T//
   xpos = 239;
   ypos = 141;
   dq_i = 85;
 
   #T//
   xpos = 240;
   ypos = 141;
   dq_i = 85;
 
   #T//
   xpos = 241;
   ypos = 141;
   dq_i = 129;
 
   #T//
   xpos = 242;
   ypos = 141;
   dq_i = 129;
 
   #T//
   xpos = 243;
   ypos = 141;
   dq_i = 164;
 
   #T//
   xpos = 244;
   ypos = 141;
   dq_i = 164;
 
   #T//
   xpos = 245;
   ypos = 141;
   dq_i = 195;
 
   #T//
   xpos = 246;
   ypos = 141;
   dq_i = 195;
 
   #T//
   xpos = 247;
   ypos = 141;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 141;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 141;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 141;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 141;
   dq_i = 106;
 
   #T//
   xpos = 252;
   ypos = 141;
   dq_i = 106;
 
   #T//
   xpos = 253;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 141;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 141;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 141;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 142;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 142;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 142;
   dq_i = 169;
 
   #T//
   xpos = 228;
   ypos = 142;
   dq_i = 169;
 
   #T//
   xpos = 229;
   ypos = 142;
   dq_i = 252;
 
   #T//
   xpos = 230;
   ypos = 142;
   dq_i = 252;
 
   #T//
   xpos = 231;
   ypos = 142;
   dq_i = 199;
 
   #T//
   xpos = 232;
   ypos = 142;
   dq_i = 199;
 
   #T//
   xpos = 233;
   ypos = 142;
   dq_i = 85;
 
   #T//
   xpos = 234;
   ypos = 142;
   dq_i = 85;
 
   #T//
   xpos = 235;
   ypos = 142;
   dq_i = 85;
 
   #T//
   xpos = 236;
   ypos = 142;
   dq_i = 85;
 
   #T//
   xpos = 237;
   ypos = 142;
   dq_i = 85;
 
   #T//
   xpos = 238;
   ypos = 142;
   dq_i = 85;
 
   #T//
   xpos = 239;
   ypos = 142;
   dq_i = 85;
 
   #T//
   xpos = 240;
   ypos = 142;
   dq_i = 85;
 
   #T//
   xpos = 241;
   ypos = 142;
   dq_i = 129;
 
   #T//
   xpos = 242;
   ypos = 142;
   dq_i = 129;
 
   #T//
   xpos = 243;
   ypos = 142;
   dq_i = 164;
 
   #T//
   xpos = 244;
   ypos = 142;
   dq_i = 164;
 
   #T//
   xpos = 245;
   ypos = 142;
   dq_i = 195;
 
   #T//
   xpos = 246;
   ypos = 142;
   dq_i = 195;
 
   #T//
   xpos = 247;
   ypos = 142;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 142;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 142;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 142;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 142;
   dq_i = 106;
 
   #T//
   xpos = 252;
   ypos = 142;
   dq_i = 106;
 
   #T//
   xpos = 253;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 142;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 142;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 142;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 143;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 143;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 143;
   dq_i = 41;
 
   #T//
   xpos = 228;
   ypos = 143;
   dq_i = 41;
 
   #T//
   xpos = 229;
   ypos = 143;
   dq_i = 170;
 
   #T//
   xpos = 230;
   ypos = 143;
   dq_i = 170;
 
   #T//
   xpos = 231;
   ypos = 143;
   dq_i = 245;
 
   #T//
   xpos = 232;
   ypos = 143;
   dq_i = 245;
 
   #T//
   xpos = 233;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 234;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 235;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 236;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 237;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 238;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 239;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 240;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 241;
   ypos = 143;
   dq_i = 232;
 
   #T//
   xpos = 242;
   ypos = 143;
   dq_i = 232;
 
   #T//
   xpos = 243;
   ypos = 143;
   dq_i = 231;
 
   #T//
   xpos = 244;
   ypos = 143;
   dq_i = 231;
 
   #T//
   xpos = 245;
   ypos = 143;
   dq_i = 251;
 
   #T//
   xpos = 246;
   ypos = 143;
   dq_i = 251;
 
   #T//
   xpos = 247;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 143;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 143;
   dq_i = 9;
 
   #T//
   xpos = 252;
   ypos = 143;
   dq_i = 9;
 
   #T//
   xpos = 253;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 143;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 143;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 143;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 144;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 144;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 144;
   dq_i = 41;
 
   #T//
   xpos = 228;
   ypos = 144;
   dq_i = 41;
 
   #T//
   xpos = 229;
   ypos = 144;
   dq_i = 170;
 
   #T//
   xpos = 230;
   ypos = 144;
   dq_i = 170;
 
   #T//
   xpos = 231;
   ypos = 144;
   dq_i = 245;
 
   #T//
   xpos = 232;
   ypos = 144;
   dq_i = 245;
 
   #T//
   xpos = 233;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 234;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 235;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 236;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 237;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 238;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 239;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 240;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 241;
   ypos = 144;
   dq_i = 232;
 
   #T//
   xpos = 242;
   ypos = 144;
   dq_i = 232;
 
   #T//
   xpos = 243;
   ypos = 144;
   dq_i = 231;
 
   #T//
   xpos = 244;
   ypos = 144;
   dq_i = 231;
 
   #T//
   xpos = 245;
   ypos = 144;
   dq_i = 251;
 
   #T//
   xpos = 246;
   ypos = 144;
   dq_i = 251;
 
   #T//
   xpos = 247;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 144;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 144;
   dq_i = 9;
 
   #T//
   xpos = 252;
   ypos = 144;
   dq_i = 9;
 
   #T//
   xpos = 253;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 144;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 144;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 144;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 145;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 145;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 145;
   dq_i = 49;
 
   #T//
   xpos = 232;
   ypos = 145;
   dq_i = 49;
 
   #T//
   xpos = 233;
   ypos = 145;
   dq_i = 84;
 
   #T//
   xpos = 234;
   ypos = 145;
   dq_i = 84;
 
   #T//
   xpos = 235;
   ypos = 145;
   dq_i = 84;
 
   #T//
   xpos = 236;
   ypos = 145;
   dq_i = 84;
 
   #T//
   xpos = 237;
   ypos = 145;
   dq_i = 84;
 
   #T//
   xpos = 238;
   ypos = 145;
   dq_i = 84;
 
   #T//
   xpos = 239;
   ypos = 145;
   dq_i = 84;
 
   #T//
   xpos = 240;
   ypos = 145;
   dq_i = 84;
 
   #T//
   xpos = 241;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 145;
   dq_i = 161;
 
   #T//
   xpos = 246;
   ypos = 145;
   dq_i = 161;
 
   #T//
   xpos = 247;
   ypos = 145;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 145;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 145;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 145;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 145;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 145;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 145;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 146;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 146;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 146;
   dq_i = 49;
 
   #T//
   xpos = 232;
   ypos = 146;
   dq_i = 49;
 
   #T//
   xpos = 233;
   ypos = 146;
   dq_i = 84;
 
   #T//
   xpos = 234;
   ypos = 146;
   dq_i = 84;
 
   #T//
   xpos = 235;
   ypos = 146;
   dq_i = 84;
 
   #T//
   xpos = 236;
   ypos = 146;
   dq_i = 84;
 
   #T//
   xpos = 237;
   ypos = 146;
   dq_i = 84;
 
   #T//
   xpos = 238;
   ypos = 146;
   dq_i = 84;
 
   #T//
   xpos = 239;
   ypos = 146;
   dq_i = 84;
 
   #T//
   xpos = 240;
   ypos = 146;
   dq_i = 84;
 
   #T//
   xpos = 241;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 146;
   dq_i = 161;
 
   #T//
   xpos = 246;
   ypos = 146;
   dq_i = 161;
 
   #T//
   xpos = 247;
   ypos = 146;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 146;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 146;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 146;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 146;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 146;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 146;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 147;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 147;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 147;
   dq_i = 127;
 
   #T//
   xpos = 246;
   ypos = 147;
   dq_i = 127;
 
   #T//
   xpos = 247;
   ypos = 147;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 147;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 147;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 147;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 147;
   dq_i = 45;
 
   #T//
   xpos = 252;
   ypos = 147;
   dq_i = 45;
 
   #T//
   xpos = 253;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 147;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 147;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 147;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 148;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 148;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 148;
   dq_i = 127;
 
   #T//
   xpos = 246;
   ypos = 148;
   dq_i = 127;
 
   #T//
   xpos = 247;
   ypos = 148;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 148;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 148;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 148;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 148;
   dq_i = 45;
 
   #T//
   xpos = 252;
   ypos = 148;
   dq_i = 45;
 
   #T//
   xpos = 253;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 148;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 148;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 148;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 149;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 149;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 149;
   dq_i = 128;
 
   #T//
   xpos = 246;
   ypos = 149;
   dq_i = 128;
 
   #T//
   xpos = 247;
   ypos = 149;
   dq_i = 253;
 
   #T//
   xpos = 248;
   ypos = 149;
   dq_i = 253;
 
   #T//
   xpos = 249;
   ypos = 149;
   dq_i = 253;
 
   #T//
   xpos = 250;
   ypos = 149;
   dq_i = 253;
 
   #T//
   xpos = 251;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 149;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 149;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 149;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 150;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 150;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 150;
   dq_i = 128;
 
   #T//
   xpos = 246;
   ypos = 150;
   dq_i = 128;
 
   #T//
   xpos = 247;
   ypos = 150;
   dq_i = 253;
 
   #T//
   xpos = 248;
   ypos = 150;
   dq_i = 253;
 
   #T//
   xpos = 249;
   ypos = 150;
   dq_i = 253;
 
   #T//
   xpos = 250;
   ypos = 150;
   dq_i = 253;
 
   #T//
   xpos = 251;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 150;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 150;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 150;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 151;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 151;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 151;
   dq_i = 127;
 
   #T//
   xpos = 246;
   ypos = 151;
   dq_i = 127;
 
   #T//
   xpos = 247;
   ypos = 151;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 151;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 151;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 151;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 151;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 151;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 151;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 152;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 152;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 152;
   dq_i = 127;
 
   #T//
   xpos = 246;
   ypos = 152;
   dq_i = 127;
 
   #T//
   xpos = 247;
   ypos = 152;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 152;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 152;
   dq_i = 252;
 
   #T//
   xpos = 250;
   ypos = 152;
   dq_i = 252;
 
   #T//
   xpos = 251;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 152;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 152;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 152;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 153;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 153;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 153;
   dq_i = 135;
 
   #T//
   xpos = 246;
   ypos = 153;
   dq_i = 135;
 
   #T//
   xpos = 247;
   ypos = 153;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 153;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 153;
   dq_i = 244;
 
   #T//
   xpos = 250;
   ypos = 153;
   dq_i = 244;
 
   #T//
   xpos = 251;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 153;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 153;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 153;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 154;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 154;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 154;
   dq_i = 135;
 
   #T//
   xpos = 246;
   ypos = 154;
   dq_i = 135;
 
   #T//
   xpos = 247;
   ypos = 154;
   dq_i = 252;
 
   #T//
   xpos = 248;
   ypos = 154;
   dq_i = 252;
 
   #T//
   xpos = 249;
   ypos = 154;
   dq_i = 244;
 
   #T//
   xpos = 250;
   ypos = 154;
   dq_i = 244;
 
   #T//
   xpos = 251;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 154;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 154;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 154;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 155;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 155;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 155;
   dq_i = 232;
 
   #T//
   xpos = 246;
   ypos = 155;
   dq_i = 232;
 
   #T//
   xpos = 247;
   ypos = 155;
   dq_i = 236;
 
   #T//
   xpos = 248;
   ypos = 155;
   dq_i = 236;
 
   #T//
   xpos = 249;
   ypos = 155;
   dq_i = 111;
 
   #T//
   xpos = 250;
   ypos = 155;
   dq_i = 111;
 
   #T//
   xpos = 251;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 155;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 155;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 155;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 156;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 156;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 156;
   dq_i = 232;
 
   #T//
   xpos = 246;
   ypos = 156;
   dq_i = 232;
 
   #T//
   xpos = 247;
   ypos = 156;
   dq_i = 236;
 
   #T//
   xpos = 248;
   ypos = 156;
   dq_i = 236;
 
   #T//
   xpos = 249;
   ypos = 156;
   dq_i = 111;
 
   #T//
   xpos = 250;
   ypos = 156;
   dq_i = 111;
 
   #T//
   xpos = 251;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 156;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 156;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 156;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 157;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 157;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 157;
   dq_i = 179;
 
   #T//
   xpos = 246;
   ypos = 157;
   dq_i = 179;
 
   #T//
   xpos = 247;
   ypos = 157;
   dq_i = 66;
 
   #T//
   xpos = 248;
   ypos = 157;
   dq_i = 66;
 
   #T//
   xpos = 249;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 157;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 157;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 157;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 158;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 158;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 158;
   dq_i = 179;
 
   #T//
   xpos = 246;
   ypos = 158;
   dq_i = 179;
 
   #T//
   xpos = 247;
   ypos = 158;
   dq_i = 66;
 
   #T//
   xpos = 248;
   ypos = 158;
   dq_i = 66;
 
   #T//
   xpos = 249;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 158;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 158;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 158;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 159;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 159;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 159;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 159;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 159;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 160;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 160;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 160;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 160;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 160;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 161;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 161;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 161;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 161;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 161;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 162;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 162;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 268;
   ypos = 162;
   dq_i = 0;
 
   #T//
   xpos = 269;
   ypos = 162;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 162;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 163;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 163;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 163;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 163;
   dq_i = 0
;
 
   #T//
   xpos = 268;
   ypos = 163;
   dq_i = 0
;
 
   #T//
   xpos = 269;
   ypos = 163;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 163;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 164;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 164;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 214;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 215;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 216;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 217;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 218;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 219;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 220;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 221;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 222;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 223;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 224;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 225;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 226;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 227;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 228;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 229;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 230;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 231;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 232;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 233;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 234;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 235;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 236;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 237;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 238;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 239;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 240;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 241;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 242;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 243;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 244;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 245;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 246;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 247;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 248;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 249;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 250;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 251;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 252;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 253;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 254;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 255;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 256;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 257;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 258;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 259;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 260;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 261;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 262;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 263;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 264;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 265;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 266;
   ypos = 164;
   dq_i = 0;
 
   #T//
   xpos = 267;
   ypos = 164;
   dq_i = 0
;
 
   #T//
   xpos = 268;
   ypos = 164;
   dq_i = 0
;
 
   #T//
   xpos = 269;
   ypos = 164;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 164;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 214;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 215;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 216;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 217;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 218;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 219;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 220;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 221;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 222;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 223;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 224;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 225;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 226;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 227;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 228;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 229;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 230;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 231;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 232;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 233;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 234;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 235;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 236;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 237;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 238;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 239;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 240;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 241;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 242;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 243;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 244;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 245;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 246;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 247;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 248;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 249;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 250;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 251;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 252;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 253;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 254;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 255;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 256;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 257;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 258;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 259;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 260;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 261;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 262;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 263;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 264;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 265;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 266;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 267;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 268;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 269;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 165;
   dq_i = 8'd0;
 
   #T//
   xpos = 211;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 212;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 213;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 214;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 215;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 216;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 217;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 218;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 219;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 220;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 221;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 222;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 223;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 224;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 225;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 226;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 227;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 228;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 229;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 230;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 231;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 232;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 233;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 234;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 235;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 236;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 237;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 238;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 239;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 240;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 241;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 242;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 243;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 244;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 245;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 246;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 247;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 248;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 249;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 250;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 251;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 252;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 253;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 254;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 255;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 256;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 257;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 258;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 259;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 260;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 261;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 262;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 263;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 264;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 265;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 266;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 267;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 268;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 269;
   ypos = 166;
   dq_i = 8'd0;
 
   #T//
   xpos = 270;
   ypos = 166;
   dq_i = 8'd0;
 
// ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** ** *
   #(T*3) //3 end 
// 80.0 ns
   rst_n      =1'b0;
end
 
always #(T/2) clk = ~clk;
 
digital_recognition u_digital_recognition(
 .clk (clk),
 .rst_n (rst_n),
 
//*binarization intgerface
 .dq_i (dq_i),
 .xpos (xpos),
 .ypos (ypos),
 .digit (digit)
);
 
 
 
endmodule
