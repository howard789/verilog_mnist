module digital_recognition #(
	parameter	[10:0]		UP			=	108,
	parameter	[10:0]		DOWN		=	164,
	parameter	[10:0]		LEFT		=	212,
	parameter	[10:0]		RIGHT		=	269,
	parameter	[10:0]		EACH_WIDE	=   2,
	parameter           	DEBIT       =   22

)(
	//system signals
	input								clk, 
	input								rst_n,
	
	//binarization 
	input			   [ 7:0]			dq_i,
	input			   [10:0]      		xpos,
	input			   [10:0]      		ypos,

	output	  reg      [ 4:0]		    digit

);

wire res_done_x784;

reg 	[ 2:0]	  done_all_res;

reg  signed [DEBIT:0]  res_0_sum;
reg  signed [DEBIT:0]  res_1_sum;
reg  signed [DEBIT:0]  res_2_sum;
reg  signed [DEBIT:0]  res_3_sum;
reg  signed [DEBIT:0]  res_4_sum;
reg  signed [DEBIT:0]  res_5_sum;
reg  signed [DEBIT:0]  res_6_sum;
reg  signed [DEBIT:0]  res_7_sum;
reg  signed [DEBIT:0]  res_8_sum;
reg  signed [DEBIT:0]  res_9_sum;



//****************************    B输入    *******************************

localparam signed [DEBIT:0]  B_0 = - 23'd4599;
localparam signed [DEBIT:0]  B_1 = - 23'd3332;
localparam signed [DEBIT:0]  B_2 = - 23'd4722;
localparam signed [DEBIT:0]  B_3 = - 23'd5087;
localparam signed [DEBIT:0]  B_4 = - 23'd3820;
localparam signed [DEBIT:0]  B_5 = - 23'd3477;
localparam signed [DEBIT:0]  B_6 = - 23'd4286;
localparam signed [DEBIT:0]  B_7 = - 23'd3446;
localparam signed [DEBIT:0]  B_8 = - 23'd7252;
localparam signed [DEBIT:0]  B_9 = - 23'd5047;


assign rst_valid =((xpos == LEFT - 1) && (ypos == UP +1)) || !rst_n;

always @ (posedge clk or negedge rst_n) begin
	if(rst_n == 1'b0) done_all_res <= 1'b0;
    else done_all_res <= {done_all_res[1:0], res_done_x784};
end

wire		  add_b;
wire		  decide_number;





always @ (posedge clk) begin
	if(!rst_n) 
		digit <= 1'b0;
		
	if(done_all_res[2]) begin	
	/*
		$monitor ($time, ,"res_0_sum = %d",res_0_sum);
		$monitor ($time, ,"res_1_sum = %d",res_1_sum);
		$monitor ($time, ,"res_2_sum = %d",res_2_sum);
		$monitor ($time, ,"res_3_sum = %d",res_3_sum);
		$monitor ($time, ,"res_4_sum = %d",res_4_sum);
		$monitor ($time, ,"res_5_sum = %d",res_5_sum);
		$monitor ($time, ,"res_6_sum = %d",res_6_sum);
		$monitor ($time, ,"res_7_sum = %d",res_7_sum);
		$monitor ($time, ,"res_8_sum = %d",res_8_sum);
		$monitor ($time, ,"res_9_sum = %d",res_9_sum);
*/
        if ((res_0_sum > res_1_sum ) &&(res_0_sum > res_2_sum ) && (res_0_sum > res_3_sum ) && (res_0_sum > res_4_sum ) && (res_0_sum > res_5_sum ) && (res_0_sum > res_6_sum ) && (res_0_sum > res_7_sum ) && (res_0_sum > res_8_sum ) && (res_0_sum > res_9_sum ) )
        	digit <= 4'd0;
		else if ((res_1_sum > res_0_sum ) &&(res_1_sum > res_2_sum ) &&(res_1_sum > res_3_sum ) &&(res_1_sum > res_4_sum ) &&(res_1_sum > res_5_sum ) &&(res_1_sum > res_6_sum ) &&(res_1_sum > res_7_sum ) &&(res_1_sum > res_8_sum ) &&(res_1_sum > res_9_sum ) )
			digit <= 4'd1;
		else if ((res_2_sum > res_0_sum ) &&(res_2_sum > res_1_sum ) &&(res_2_sum > res_3_sum ) &&(res_2_sum > res_4_sum ) &&(res_2_sum > res_5_sum ) &&(res_2_sum > res_6_sum ) &&(res_2_sum > res_7_sum ) &&(res_2_sum > res_8_sum ) &&(res_2_sum > res_9_sum ) )
     		digit <= 4'd2;
     	else if ((res_3_sum > res_0_sum ) &&(res_3_sum > res_1_sum ) &&(res_3_sum > res_2_sum ) &&(res_3_sum > res_4_sum ) &&(res_3_sum > res_5_sum ) &&(res_3_sum > res_6_sum ) &&(res_3_sum > res_7_sum ) &&(res_3_sum > res_8_sum ) &&(res_3_sum > res_9_sum ) )
		     digit <= 4'd3;
		else if ((res_4_sum > res_0_sum ) &&(res_4_sum > res_1_sum ) &&(res_4_sum > res_2_sum ) &&(res_4_sum > res_3_sum ) &&(res_4_sum > res_5_sum ) &&(res_4_sum > res_6_sum ) &&(res_4_sum > res_7_sum ) &&(res_4_sum > res_8_sum ) &&(res_4_sum > res_9_sum ) )
		     digit <= 4'd4;
		else if ((res_5_sum > res_0_sum ) &&(res_5_sum > res_1_sum ) &&(res_5_sum > res_2_sum ) &&(res_5_sum > res_3_sum ) &&(res_5_sum > res_4_sum ) &&(res_5_sum > res_6_sum ) &&(res_5_sum > res_7_sum ) &&(res_5_sum > res_8_sum ) &&(res_5_sum > res_9_sum ) )
		     digit <= 4'd5;
		else if ((res_6_sum > res_0_sum ) &&(res_6_sum > res_1_sum ) &&(res_6_sum > res_2_sum ) &&(res_6_sum > res_3_sum ) &&(res_6_sum > res_4_sum ) &&(res_6_sum > res_5_sum ) &&(res_6_sum > res_7_sum ) &&(res_6_sum > res_8_sum ) &&(res_6_sum > res_9_sum ) )
		     digit <= 4'd6;
		else if ((res_7_sum > res_0_sum ) &&(res_7_sum > res_1_sum ) &&(res_7_sum > res_2_sum ) &&(res_7_sum > res_3_sum ) &&(res_7_sum > res_4_sum ) &&(res_7_sum > res_5_sum ) &&(res_7_sum > res_6_sum ) &&(res_7_sum > res_8_sum ) &&(res_7_sum > res_9_sum ) )
		     digit <= 4'd7;
		else if ((res_8_sum > res_0_sum ) &&(res_8_sum > res_1_sum ) &&(res_8_sum > res_2_sum ) &&(res_8_sum > res_3_sum ) &&(res_8_sum > res_4_sum ) &&(res_8_sum > res_5_sum ) &&(res_8_sum > res_6_sum ) &&(res_8_sum > res_7_sum ) &&(res_8_sum > res_9_sum ) )
		     digit <= 4'd8;
		else if ((res_9_sum > res_0_sum ) &&(res_9_sum > res_1_sum ) &&(res_9_sum > res_2_sum ) &&(res_9_sum > res_3_sum ) &&(res_9_sum > res_4_sum ) &&(res_9_sum > res_5_sum ) &&(res_9_sum > res_6_sum ) &&(res_9_sum > res_7_sum ) &&(res_9_sum > res_8_sum ) )
		     digit <= 4'd9;
		else 
			digit <= 4'd10;     

    end 
end

//****************************    wire    *******************************
wire res_done_x1;
wire res_done_x2;
wire res_done_x3;
wire res_done_x4;
wire res_done_x5;
wire res_done_x6;
wire res_done_x7;
wire res_done_x8;
wire res_done_x9;
wire res_done_x10;
wire res_done_x11;
wire res_done_x12;
wire res_done_x13;
wire res_done_x14;
wire res_done_x15;
wire res_done_x16;
wire res_done_x17;
wire res_done_x18;
wire res_done_x19;
wire res_done_x20;
wire res_done_x21;
wire res_done_x22;
wire res_done_x23;
wire res_done_x24;
wire res_done_x25;
wire res_done_x26;
wire res_done_x27;
wire res_done_x28;
wire res_done_x29;
wire res_done_x30;
wire res_done_x31;
wire res_done_x32;
wire res_done_x33;
wire res_done_x34;
wire res_done_x35;
wire res_done_x36;
wire res_done_x37;
wire res_done_x38;
wire res_done_x39;
wire res_done_x40;
wire res_done_x41;
wire res_done_x42;
wire res_done_x43;
wire res_done_x44;
wire res_done_x45;
wire res_done_x46;
wire res_done_x47;
wire res_done_x48;
wire res_done_x49;
wire res_done_x50;
wire res_done_x51;
wire res_done_x52;
wire res_done_x53;
wire res_done_x54;
wire res_done_x55;
wire res_done_x56;
wire res_done_x57;
wire res_done_x58;
wire res_done_x59;
wire res_done_x60;
wire res_done_x61;
wire res_done_x62;
wire res_done_x63;
wire res_done_x64;
wire res_done_x65;
wire res_done_x66;
wire res_done_x67;
wire res_done_x68;
wire res_done_x69;
wire res_done_x70;
wire res_done_x71;
wire res_done_x72;
wire res_done_x73;
wire res_done_x74;
wire res_done_x75;
wire res_done_x76;
wire res_done_x77;
wire res_done_x78;
wire res_done_x79;
wire res_done_x80;
wire res_done_x81;
wire res_done_x82;
wire res_done_x83;
wire res_done_x84;
wire res_done_x85;
wire res_done_x86;
wire res_done_x87;
wire res_done_x88;
wire res_done_x89;
wire res_done_x90;
wire res_done_x91;
wire res_done_x92;
wire res_done_x93;
wire res_done_x94;
wire res_done_x95;
wire res_done_x96;
wire res_done_x97;
wire res_done_x98;
wire res_done_x99;
wire res_done_x100;
wire res_done_x101;
wire res_done_x102;
wire res_done_x103;
wire res_done_x104;
wire res_done_x105;
wire res_done_x106;
wire res_done_x107;
wire res_done_x108;
wire res_done_x109;
wire res_done_x110;
wire res_done_x111;
wire res_done_x112;
wire res_done_x113;
wire res_done_x114;
wire res_done_x115;
wire res_done_x116;
wire res_done_x117;
wire res_done_x118;
wire res_done_x119;
wire res_done_x120;
wire res_done_x121;
wire res_done_x122;
wire res_done_x123;
wire res_done_x124;
wire res_done_x125;
wire res_done_x126;
wire res_done_x127;
wire res_done_x128;
wire res_done_x129;
wire res_done_x130;
wire res_done_x131;
wire res_done_x132;
wire res_done_x133;
wire res_done_x134;
wire res_done_x135;
wire res_done_x136;
wire res_done_x137;
wire res_done_x138;
wire res_done_x139;
wire res_done_x140;
wire res_done_x141;
wire res_done_x142;
wire res_done_x143;
wire res_done_x144;
wire res_done_x145;
wire res_done_x146;
wire res_done_x147;
wire res_done_x148;
wire res_done_x149;
wire res_done_x150;
wire res_done_x151;
wire res_done_x152;
wire res_done_x153;
wire res_done_x154;
wire res_done_x155;
wire res_done_x156;
wire res_done_x157;
wire res_done_x158;
wire res_done_x159;
wire res_done_x160;
wire res_done_x161;
wire res_done_x162;
wire res_done_x163;
wire res_done_x164;
wire res_done_x165;
wire res_done_x166;
wire res_done_x167;
wire res_done_x168;
wire res_done_x169;
wire res_done_x170;
wire res_done_x171;
wire res_done_x172;
wire res_done_x173;
wire res_done_x174;
wire res_done_x175;
wire res_done_x176;
wire res_done_x177;
wire res_done_x178;
wire res_done_x179;
wire res_done_x180;
wire res_done_x181;
wire res_done_x182;
wire res_done_x183;
wire res_done_x184;
wire res_done_x185;
wire res_done_x186;
wire res_done_x187;
wire res_done_x188;
wire res_done_x189;
wire res_done_x190;
wire res_done_x191;
wire res_done_x192;
wire res_done_x193;
wire res_done_x194;
wire res_done_x195;
wire res_done_x196;
wire res_done_x197;
wire res_done_x198;
wire res_done_x199;
wire res_done_x200;
wire res_done_x201;
wire res_done_x202;
wire res_done_x203;
wire res_done_x204;
wire res_done_x205;
wire res_done_x206;
wire res_done_x207;
wire res_done_x208;
wire res_done_x209;
wire res_done_x210;
wire res_done_x211;
wire res_done_x212;
wire res_done_x213;
wire res_done_x214;
wire res_done_x215;
wire res_done_x216;
wire res_done_x217;
wire res_done_x218;
wire res_done_x219;
wire res_done_x220;
wire res_done_x221;
wire res_done_x222;
wire res_done_x223;
wire res_done_x224;
wire res_done_x225;
wire res_done_x226;
wire res_done_x227;
wire res_done_x228;
wire res_done_x229;
wire res_done_x230;
wire res_done_x231;
wire res_done_x232;
wire res_done_x233;
wire res_done_x234;
wire res_done_x235;
wire res_done_x236;
wire res_done_x237;
wire res_done_x238;
wire res_done_x239;
wire res_done_x240;
wire res_done_x241;
wire res_done_x242;
wire res_done_x243;
wire res_done_x244;
wire res_done_x245;
wire res_done_x246;
wire res_done_x247;
wire res_done_x248;
wire res_done_x249;
wire res_done_x250;
wire res_done_x251;
wire res_done_x252;
wire res_done_x253;
wire res_done_x254;
wire res_done_x255;
wire res_done_x256;
wire res_done_x257;
wire res_done_x258;
wire res_done_x259;
wire res_done_x260;
wire res_done_x261;
wire res_done_x262;
wire res_done_x263;
wire res_done_x264;
wire res_done_x265;
wire res_done_x266;
wire res_done_x267;
wire res_done_x268;
wire res_done_x269;
wire res_done_x270;
wire res_done_x271;
wire res_done_x272;
wire res_done_x273;
wire res_done_x274;
wire res_done_x275;
wire res_done_x276;
wire res_done_x277;
wire res_done_x278;
wire res_done_x279;
wire res_done_x280;
wire res_done_x281;
wire res_done_x282;
wire res_done_x283;
wire res_done_x284;
wire res_done_x285;
wire res_done_x286;
wire res_done_x287;
wire res_done_x288;
wire res_done_x289;
wire res_done_x290;
wire res_done_x291;
wire res_done_x292;
wire res_done_x293;
wire res_done_x294;
wire res_done_x295;
wire res_done_x296;
wire res_done_x297;
wire res_done_x298;
wire res_done_x299;
wire res_done_x300;
wire res_done_x301;
wire res_done_x302;
wire res_done_x303;
wire res_done_x304;
wire res_done_x305;
wire res_done_x306;
wire res_done_x307;
wire res_done_x308;
wire res_done_x309;
wire res_done_x310;
wire res_done_x311;
wire res_done_x312;
wire res_done_x313;
wire res_done_x314;
wire res_done_x315;
wire res_done_x316;
wire res_done_x317;
wire res_done_x318;
wire res_done_x319;
wire res_done_x320;
wire res_done_x321;
wire res_done_x322;
wire res_done_x323;
wire res_done_x324;
wire res_done_x325;
wire res_done_x326;
wire res_done_x327;
wire res_done_x328;
wire res_done_x329;
wire res_done_x330;
wire res_done_x331;
wire res_done_x332;
wire res_done_x333;
wire res_done_x334;
wire res_done_x335;
wire res_done_x336;
wire res_done_x337;
wire res_done_x338;
wire res_done_x339;
wire res_done_x340;
wire res_done_x341;
wire res_done_x342;
wire res_done_x343;
wire res_done_x344;
wire res_done_x345;
wire res_done_x346;
wire res_done_x347;
wire res_done_x348;
wire res_done_x349;
wire res_done_x350;
wire res_done_x351;
wire res_done_x352;
wire res_done_x353;
wire res_done_x354;
wire res_done_x355;
wire res_done_x356;
wire res_done_x357;
wire res_done_x358;
wire res_done_x359;
wire res_done_x360;
wire res_done_x361;
wire res_done_x362;
wire res_done_x363;
wire res_done_x364;
wire res_done_x365;
wire res_done_x366;
wire res_done_x367;
wire res_done_x368;
wire res_done_x369;
wire res_done_x370;
wire res_done_x371;
wire res_done_x372;
wire res_done_x373;
wire res_done_x374;
wire res_done_x375;
wire res_done_x376;
wire res_done_x377;
wire res_done_x378;
wire res_done_x379;
wire res_done_x380;
wire res_done_x381;
wire res_done_x382;
wire res_done_x383;
wire res_done_x384;
wire res_done_x385;
wire res_done_x386;
wire res_done_x387;
wire res_done_x388;
wire res_done_x389;
wire res_done_x390;
wire res_done_x391;
wire res_done_x392;
wire res_done_x393;
wire res_done_x394;
wire res_done_x395;
wire res_done_x396;
wire res_done_x397;
wire res_done_x398;
wire res_done_x399;
wire res_done_x400;
wire res_done_x401;
wire res_done_x402;
wire res_done_x403;
wire res_done_x404;
wire res_done_x405;
wire res_done_x406;
wire res_done_x407;
wire res_done_x408;
wire res_done_x409;
wire res_done_x410;
wire res_done_x411;
wire res_done_x412;
wire res_done_x413;
wire res_done_x414;
wire res_done_x415;
wire res_done_x416;
wire res_done_x417;
wire res_done_x418;
wire res_done_x419;
wire res_done_x420;
wire res_done_x421;
wire res_done_x422;
wire res_done_x423;
wire res_done_x424;
wire res_done_x425;
wire res_done_x426;
wire res_done_x427;
wire res_done_x428;
wire res_done_x429;
wire res_done_x430;
wire res_done_x431;
wire res_done_x432;
wire res_done_x433;
wire res_done_x434;
wire res_done_x435;
wire res_done_x436;
wire res_done_x437;
wire res_done_x438;
wire res_done_x439;
wire res_done_x440;
wire res_done_x441;
wire res_done_x442;
wire res_done_x443;
wire res_done_x444;
wire res_done_x445;
wire res_done_x446;
wire res_done_x447;
wire res_done_x448;
wire res_done_x449;
wire res_done_x450;
wire res_done_x451;
wire res_done_x452;
wire res_done_x453;
wire res_done_x454;
wire res_done_x455;
wire res_done_x456;
wire res_done_x457;
wire res_done_x458;
wire res_done_x459;
wire res_done_x460;
wire res_done_x461;
wire res_done_x462;
wire res_done_x463;
wire res_done_x464;
wire res_done_x465;
wire res_done_x466;
wire res_done_x467;
wire res_done_x468;
wire res_done_x469;
wire res_done_x470;
wire res_done_x471;
wire res_done_x472;
wire res_done_x473;
wire res_done_x474;
wire res_done_x475;
wire res_done_x476;
wire res_done_x477;
wire res_done_x478;
wire res_done_x479;
wire res_done_x480;
wire res_done_x481;
wire res_done_x482;
wire res_done_x483;
wire res_done_x484;
wire res_done_x485;
wire res_done_x486;
wire res_done_x487;
wire res_done_x488;
wire res_done_x489;
wire res_done_x490;
wire res_done_x491;
wire res_done_x492;
wire res_done_x493;
wire res_done_x494;
wire res_done_x495;
wire res_done_x496;
wire res_done_x497;
wire res_done_x498;
wire res_done_x499;
wire res_done_x500;
wire res_done_x501;
wire res_done_x502;
wire res_done_x503;
wire res_done_x504;
wire res_done_x505;
wire res_done_x506;
wire res_done_x507;
wire res_done_x508;
wire res_done_x509;
wire res_done_x510;
wire res_done_x511;
wire res_done_x512;
wire res_done_x513;
wire res_done_x514;
wire res_done_x515;
wire res_done_x516;
wire res_done_x517;
wire res_done_x518;
wire res_done_x519;
wire res_done_x520;
wire res_done_x521;
wire res_done_x522;
wire res_done_x523;
wire res_done_x524;
wire res_done_x525;
wire res_done_x526;
wire res_done_x527;
wire res_done_x528;
wire res_done_x529;
wire res_done_x530;
wire res_done_x531;
wire res_done_x532;
wire res_done_x533;
wire res_done_x534;
wire res_done_x535;
wire res_done_x536;
wire res_done_x537;
wire res_done_x538;
wire res_done_x539;
wire res_done_x540;
wire res_done_x541;
wire res_done_x542;
wire res_done_x543;
wire res_done_x544;
wire res_done_x545;
wire res_done_x546;
wire res_done_x547;
wire res_done_x548;
wire res_done_x549;
wire res_done_x550;
wire res_done_x551;
wire res_done_x552;
wire res_done_x553;
wire res_done_x554;
wire res_done_x555;
wire res_done_x556;
wire res_done_x557;
wire res_done_x558;
wire res_done_x559;
wire res_done_x560;
wire res_done_x561;
wire res_done_x562;
wire res_done_x563;
wire res_done_x564;
wire res_done_x565;
wire res_done_x566;
wire res_done_x567;
wire res_done_x568;
wire res_done_x569;
wire res_done_x570;
wire res_done_x571;
wire res_done_x572;
wire res_done_x573;
wire res_done_x574;
wire res_done_x575;
wire res_done_x576;
wire res_done_x577;
wire res_done_x578;
wire res_done_x579;
wire res_done_x580;
wire res_done_x581;
wire res_done_x582;
wire res_done_x583;
wire res_done_x584;
wire res_done_x585;
wire res_done_x586;
wire res_done_x587;
wire res_done_x588;
wire res_done_x589;
wire res_done_x590;
wire res_done_x591;
wire res_done_x592;
wire res_done_x593;
wire res_done_x594;
wire res_done_x595;
wire res_done_x596;
wire res_done_x597;
wire res_done_x598;
wire res_done_x599;
wire res_done_x600;
wire res_done_x601;
wire res_done_x602;
wire res_done_x603;
wire res_done_x604;
wire res_done_x605;
wire res_done_x606;
wire res_done_x607;
wire res_done_x608;
wire res_done_x609;
wire res_done_x610;
wire res_done_x611;
wire res_done_x612;
wire res_done_x613;
wire res_done_x614;
wire res_done_x615;
wire res_done_x616;
wire res_done_x617;
wire res_done_x618;
wire res_done_x619;
wire res_done_x620;
wire res_done_x621;
wire res_done_x622;
wire res_done_x623;
wire res_done_x624;
wire res_done_x625;
wire res_done_x626;
wire res_done_x627;
wire res_done_x628;
wire res_done_x629;
wire res_done_x630;
wire res_done_x631;
wire res_done_x632;
wire res_done_x633;
wire res_done_x634;
wire res_done_x635;
wire res_done_x636;
wire res_done_x637;
wire res_done_x638;
wire res_done_x639;
wire res_done_x640;
wire res_done_x641;
wire res_done_x642;
wire res_done_x643;
wire res_done_x644;
wire res_done_x645;
wire res_done_x646;
wire res_done_x647;
wire res_done_x648;
wire res_done_x649;
wire res_done_x650;
wire res_done_x651;
wire res_done_x652;
wire res_done_x653;
wire res_done_x654;
wire res_done_x655;
wire res_done_x656;
wire res_done_x657;
wire res_done_x658;
wire res_done_x659;
wire res_done_x660;
wire res_done_x661;
wire res_done_x662;
wire res_done_x663;
wire res_done_x664;
wire res_done_x665;
wire res_done_x666;
wire res_done_x667;
wire res_done_x668;
wire res_done_x669;
wire res_done_x670;
wire res_done_x671;
wire res_done_x672;
wire res_done_x673;
wire res_done_x674;
wire res_done_x675;
wire res_done_x676;
wire res_done_x677;
wire res_done_x678;
wire res_done_x679;
wire res_done_x680;
wire res_done_x681;
wire res_done_x682;
wire res_done_x683;
wire res_done_x684;
wire res_done_x685;
wire res_done_x686;
wire res_done_x687;
wire res_done_x688;
wire res_done_x689;
wire res_done_x690;
wire res_done_x691;
wire res_done_x692;
wire res_done_x693;
wire res_done_x694;
wire res_done_x695;
wire res_done_x696;
wire res_done_x697;
wire res_done_x698;
wire res_done_x699;
wire res_done_x700;
wire res_done_x701;
wire res_done_x702;
wire res_done_x703;
wire res_done_x704;
wire res_done_x705;
wire res_done_x706;
wire res_done_x707;
wire res_done_x708;
wire res_done_x709;
wire res_done_x710;
wire res_done_x711;
wire res_done_x712;
wire res_done_x713;
wire res_done_x714;
wire res_done_x715;
wire res_done_x716;
wire res_done_x717;
wire res_done_x718;
wire res_done_x719;
wire res_done_x720;
wire res_done_x721;
wire res_done_x722;
wire res_done_x723;
wire res_done_x724;
wire res_done_x725;
wire res_done_x726;
wire res_done_x727;
wire res_done_x728;
wire res_done_x729;
wire res_done_x730;
wire res_done_x731;
wire res_done_x732;
wire res_done_x733;
wire res_done_x734;
wire res_done_x735;
wire res_done_x736;
wire res_done_x737;
wire res_done_x738;
wire res_done_x739;
wire res_done_x740;
wire res_done_x741;
wire res_done_x742;
wire res_done_x743;
wire res_done_x744;
wire res_done_x745;
wire res_done_x746;
wire res_done_x747;
wire res_done_x748;
wire res_done_x749;
wire res_done_x750;
wire res_done_x751;
wire res_done_x752;
wire res_done_x753;
wire res_done_x754;
wire res_done_x755;
wire res_done_x756;
wire res_done_x757;
wire res_done_x758;
wire res_done_x759;
wire res_done_x760;
wire res_done_x761;
wire res_done_x762;
wire res_done_x763;
wire res_done_x764;
wire res_done_x765;
wire res_done_x766;
wire res_done_x767;
wire res_done_x768;
wire res_done_x769;
wire res_done_x770;
wire res_done_x771;
wire res_done_x772;
wire res_done_x773;
wire res_done_x774;
wire res_done_x775;
wire res_done_x776;
wire res_done_x777;
wire res_done_x778;
wire res_done_x779;
wire res_done_x780;
wire res_done_x781;
wire res_done_x782;
wire res_done_x783;
// wire res_done_x784;


wire signed [DEBIT:0] score_0_x1;
wire signed [DEBIT:0] score_0_x2;
wire signed [DEBIT:0] score_0_x3;
wire signed [DEBIT:0] score_0_x4;
wire signed [DEBIT:0] score_0_x5;
wire signed [DEBIT:0] score_0_x6;
wire signed [DEBIT:0] score_0_x7;
wire signed [DEBIT:0] score_0_x8;
wire signed [DEBIT:0] score_0_x9;
wire signed [DEBIT:0] score_0_x10;
wire signed [DEBIT:0] score_0_x11;
wire signed [DEBIT:0] score_0_x12;
wire signed [DEBIT:0] score_0_x13;
wire signed [DEBIT:0] score_0_x14;
wire signed [DEBIT:0] score_0_x15;
wire signed [DEBIT:0] score_0_x16;
wire signed [DEBIT:0] score_0_x17;
wire signed [DEBIT:0] score_0_x18;
wire signed [DEBIT:0] score_0_x19;
wire signed [DEBIT:0] score_0_x20;
wire signed [DEBIT:0] score_0_x21;
wire signed [DEBIT:0] score_0_x22;
wire signed [DEBIT:0] score_0_x23;
wire signed [DEBIT:0] score_0_x24;
wire signed [DEBIT:0] score_0_x25;
wire signed [DEBIT:0] score_0_x26;
wire signed [DEBIT:0] score_0_x27;
wire signed [DEBIT:0] score_0_x28;
wire signed [DEBIT:0] score_0_x29;
wire signed [DEBIT:0] score_0_x30;
wire signed [DEBIT:0] score_0_x31;
wire signed [DEBIT:0] score_0_x32;
wire signed [DEBIT:0] score_0_x33;
wire signed [DEBIT:0] score_0_x34;
wire signed [DEBIT:0] score_0_x35;
wire signed [DEBIT:0] score_0_x36;
wire signed [DEBIT:0] score_0_x37;
wire signed [DEBIT:0] score_0_x38;
wire signed [DEBIT:0] score_0_x39;
wire signed [DEBIT:0] score_0_x40;
wire signed [DEBIT:0] score_0_x41;
wire signed [DEBIT:0] score_0_x42;
wire signed [DEBIT:0] score_0_x43;
wire signed [DEBIT:0] score_0_x44;
wire signed [DEBIT:0] score_0_x45;
wire signed [DEBIT:0] score_0_x46;
wire signed [DEBIT:0] score_0_x47;
wire signed [DEBIT:0] score_0_x48;
wire signed [DEBIT:0] score_0_x49;
wire signed [DEBIT:0] score_0_x50;
wire signed [DEBIT:0] score_0_x51;
wire signed [DEBIT:0] score_0_x52;
wire signed [DEBIT:0] score_0_x53;
wire signed [DEBIT:0] score_0_x54;
wire signed [DEBIT:0] score_0_x55;
wire signed [DEBIT:0] score_0_x56;
wire signed [DEBIT:0] score_0_x57;
wire signed [DEBIT:0] score_0_x58;
wire signed [DEBIT:0] score_0_x59;
wire signed [DEBIT:0] score_0_x60;
wire signed [DEBIT:0] score_0_x61;
wire signed [DEBIT:0] score_0_x62;
wire signed [DEBIT:0] score_0_x63;
wire signed [DEBIT:0] score_0_x64;
wire signed [DEBIT:0] score_0_x65;
wire signed [DEBIT:0] score_0_x66;
wire signed [DEBIT:0] score_0_x67;
wire signed [DEBIT:0] score_0_x68;
wire signed [DEBIT:0] score_0_x69;
wire signed [DEBIT:0] score_0_x70;
wire signed [DEBIT:0] score_0_x71;
wire signed [DEBIT:0] score_0_x72;
wire signed [DEBIT:0] score_0_x73;
wire signed [DEBIT:0] score_0_x74;
wire signed [DEBIT:0] score_0_x75;
wire signed [DEBIT:0] score_0_x76;
wire signed [DEBIT:0] score_0_x77;
wire signed [DEBIT:0] score_0_x78;
wire signed [DEBIT:0] score_0_x79;
wire signed [DEBIT:0] score_0_x80;
wire signed [DEBIT:0] score_0_x81;
wire signed [DEBIT:0] score_0_x82;
wire signed [DEBIT:0] score_0_x83;
wire signed [DEBIT:0] score_0_x84;
wire signed [DEBIT:0] score_0_x85;
wire signed [DEBIT:0] score_0_x86;
wire signed [DEBIT:0] score_0_x87;
wire signed [DEBIT:0] score_0_x88;
wire signed [DEBIT:0] score_0_x89;
wire signed [DEBIT:0] score_0_x90;
wire signed [DEBIT:0] score_0_x91;
wire signed [DEBIT:0] score_0_x92;
wire signed [DEBIT:0] score_0_x93;
wire signed [DEBIT:0] score_0_x94;
wire signed [DEBIT:0] score_0_x95;
wire signed [DEBIT:0] score_0_x96;
wire signed [DEBIT:0] score_0_x97;
wire signed [DEBIT:0] score_0_x98;
wire signed [DEBIT:0] score_0_x99;
wire signed [DEBIT:0] score_0_x100;
wire signed [DEBIT:0] score_0_x101;
wire signed [DEBIT:0] score_0_x102;
wire signed [DEBIT:0] score_0_x103;
wire signed [DEBIT:0] score_0_x104;
wire signed [DEBIT:0] score_0_x105;
wire signed [DEBIT:0] score_0_x106;
wire signed [DEBIT:0] score_0_x107;
wire signed [DEBIT:0] score_0_x108;
wire signed [DEBIT:0] score_0_x109;
wire signed [DEBIT:0] score_0_x110;
wire signed [DEBIT:0] score_0_x111;
wire signed [DEBIT:0] score_0_x112;
wire signed [DEBIT:0] score_0_x113;
wire signed [DEBIT:0] score_0_x114;
wire signed [DEBIT:0] score_0_x115;
wire signed [DEBIT:0] score_0_x116;
wire signed [DEBIT:0] score_0_x117;
wire signed [DEBIT:0] score_0_x118;
wire signed [DEBIT:0] score_0_x119;
wire signed [DEBIT:0] score_0_x120;
wire signed [DEBIT:0] score_0_x121;
wire signed [DEBIT:0] score_0_x122;
wire signed [DEBIT:0] score_0_x123;
wire signed [DEBIT:0] score_0_x124;
wire signed [DEBIT:0] score_0_x125;
wire signed [DEBIT:0] score_0_x126;
wire signed [DEBIT:0] score_0_x127;
wire signed [DEBIT:0] score_0_x128;
wire signed [DEBIT:0] score_0_x129;
wire signed [DEBIT:0] score_0_x130;
wire signed [DEBIT:0] score_0_x131;
wire signed [DEBIT:0] score_0_x132;
wire signed [DEBIT:0] score_0_x133;
wire signed [DEBIT:0] score_0_x134;
wire signed [DEBIT:0] score_0_x135;
wire signed [DEBIT:0] score_0_x136;
wire signed [DEBIT:0] score_0_x137;
wire signed [DEBIT:0] score_0_x138;
wire signed [DEBIT:0] score_0_x139;
wire signed [DEBIT:0] score_0_x140;
wire signed [DEBIT:0] score_0_x141;
wire signed [DEBIT:0] score_0_x142;
wire signed [DEBIT:0] score_0_x143;
wire signed [DEBIT:0] score_0_x144;
wire signed [DEBIT:0] score_0_x145;
wire signed [DEBIT:0] score_0_x146;
wire signed [DEBIT:0] score_0_x147;
wire signed [DEBIT:0] score_0_x148;
wire signed [DEBIT:0] score_0_x149;
wire signed [DEBIT:0] score_0_x150;
wire signed [DEBIT:0] score_0_x151;
wire signed [DEBIT:0] score_0_x152;
wire signed [DEBIT:0] score_0_x153;
wire signed [DEBIT:0] score_0_x154;
wire signed [DEBIT:0] score_0_x155;
wire signed [DEBIT:0] score_0_x156;
wire signed [DEBIT:0] score_0_x157;
wire signed [DEBIT:0] score_0_x158;
wire signed [DEBIT:0] score_0_x159;
wire signed [DEBIT:0] score_0_x160;
wire signed [DEBIT:0] score_0_x161;
wire signed [DEBIT:0] score_0_x162;
wire signed [DEBIT:0] score_0_x163;
wire signed [DEBIT:0] score_0_x164;
wire signed [DEBIT:0] score_0_x165;
wire signed [DEBIT:0] score_0_x166;
wire signed [DEBIT:0] score_0_x167;
wire signed [DEBIT:0] score_0_x168;
wire signed [DEBIT:0] score_0_x169;
wire signed [DEBIT:0] score_0_x170;
wire signed [DEBIT:0] score_0_x171;
wire signed [DEBIT:0] score_0_x172;
wire signed [DEBIT:0] score_0_x173;
wire signed [DEBIT:0] score_0_x174;
wire signed [DEBIT:0] score_0_x175;
wire signed [DEBIT:0] score_0_x176;
wire signed [DEBIT:0] score_0_x177;
wire signed [DEBIT:0] score_0_x178;
wire signed [DEBIT:0] score_0_x179;
wire signed [DEBIT:0] score_0_x180;
wire signed [DEBIT:0] score_0_x181;
wire signed [DEBIT:0] score_0_x182;
wire signed [DEBIT:0] score_0_x183;
wire signed [DEBIT:0] score_0_x184;
wire signed [DEBIT:0] score_0_x185;
wire signed [DEBIT:0] score_0_x186;
wire signed [DEBIT:0] score_0_x187;
wire signed [DEBIT:0] score_0_x188;
wire signed [DEBIT:0] score_0_x189;
wire signed [DEBIT:0] score_0_x190;
wire signed [DEBIT:0] score_0_x191;
wire signed [DEBIT:0] score_0_x192;
wire signed [DEBIT:0] score_0_x193;
wire signed [DEBIT:0] score_0_x194;
wire signed [DEBIT:0] score_0_x195;
wire signed [DEBIT:0] score_0_x196;
wire signed [DEBIT:0] score_0_x197;
wire signed [DEBIT:0] score_0_x198;
wire signed [DEBIT:0] score_0_x199;
wire signed [DEBIT:0] score_0_x200;
wire signed [DEBIT:0] score_0_x201;
wire signed [DEBIT:0] score_0_x202;
wire signed [DEBIT:0] score_0_x203;
wire signed [DEBIT:0] score_0_x204;
wire signed [DEBIT:0] score_0_x205;
wire signed [DEBIT:0] score_0_x206;
wire signed [DEBIT:0] score_0_x207;
wire signed [DEBIT:0] score_0_x208;
wire signed [DEBIT:0] score_0_x209;
wire signed [DEBIT:0] score_0_x210;
wire signed [DEBIT:0] score_0_x211;
wire signed [DEBIT:0] score_0_x212;
wire signed [DEBIT:0] score_0_x213;
wire signed [DEBIT:0] score_0_x214;
wire signed [DEBIT:0] score_0_x215;
wire signed [DEBIT:0] score_0_x216;
wire signed [DEBIT:0] score_0_x217;
wire signed [DEBIT:0] score_0_x218;
wire signed [DEBIT:0] score_0_x219;
wire signed [DEBIT:0] score_0_x220;
wire signed [DEBIT:0] score_0_x221;
wire signed [DEBIT:0] score_0_x222;
wire signed [DEBIT:0] score_0_x223;
wire signed [DEBIT:0] score_0_x224;
wire signed [DEBIT:0] score_0_x225;
wire signed [DEBIT:0] score_0_x226;
wire signed [DEBIT:0] score_0_x227;
wire signed [DEBIT:0] score_0_x228;
wire signed [DEBIT:0] score_0_x229;
wire signed [DEBIT:0] score_0_x230;
wire signed [DEBIT:0] score_0_x231;
wire signed [DEBIT:0] score_0_x232;
wire signed [DEBIT:0] score_0_x233;
wire signed [DEBIT:0] score_0_x234;
wire signed [DEBIT:0] score_0_x235;
wire signed [DEBIT:0] score_0_x236;
wire signed [DEBIT:0] score_0_x237;
wire signed [DEBIT:0] score_0_x238;
wire signed [DEBIT:0] score_0_x239;
wire signed [DEBIT:0] score_0_x240;
wire signed [DEBIT:0] score_0_x241;
wire signed [DEBIT:0] score_0_x242;
wire signed [DEBIT:0] score_0_x243;
wire signed [DEBIT:0] score_0_x244;
wire signed [DEBIT:0] score_0_x245;
wire signed [DEBIT:0] score_0_x246;
wire signed [DEBIT:0] score_0_x247;
wire signed [DEBIT:0] score_0_x248;
wire signed [DEBIT:0] score_0_x249;
wire signed [DEBIT:0] score_0_x250;
wire signed [DEBIT:0] score_0_x251;
wire signed [DEBIT:0] score_0_x252;
wire signed [DEBIT:0] score_0_x253;
wire signed [DEBIT:0] score_0_x254;
wire signed [DEBIT:0] score_0_x255;
wire signed [DEBIT:0] score_0_x256;
wire signed [DEBIT:0] score_0_x257;
wire signed [DEBIT:0] score_0_x258;
wire signed [DEBIT:0] score_0_x259;
wire signed [DEBIT:0] score_0_x260;
wire signed [DEBIT:0] score_0_x261;
wire signed [DEBIT:0] score_0_x262;
wire signed [DEBIT:0] score_0_x263;
wire signed [DEBIT:0] score_0_x264;
wire signed [DEBIT:0] score_0_x265;
wire signed [DEBIT:0] score_0_x266;
wire signed [DEBIT:0] score_0_x267;
wire signed [DEBIT:0] score_0_x268;
wire signed [DEBIT:0] score_0_x269;
wire signed [DEBIT:0] score_0_x270;
wire signed [DEBIT:0] score_0_x271;
wire signed [DEBIT:0] score_0_x272;
wire signed [DEBIT:0] score_0_x273;
wire signed [DEBIT:0] score_0_x274;
wire signed [DEBIT:0] score_0_x275;
wire signed [DEBIT:0] score_0_x276;
wire signed [DEBIT:0] score_0_x277;
wire signed [DEBIT:0] score_0_x278;
wire signed [DEBIT:0] score_0_x279;
wire signed [DEBIT:0] score_0_x280;
wire signed [DEBIT:0] score_0_x281;
wire signed [DEBIT:0] score_0_x282;
wire signed [DEBIT:0] score_0_x283;
wire signed [DEBIT:0] score_0_x284;
wire signed [DEBIT:0] score_0_x285;
wire signed [DEBIT:0] score_0_x286;
wire signed [DEBIT:0] score_0_x287;
wire signed [DEBIT:0] score_0_x288;
wire signed [DEBIT:0] score_0_x289;
wire signed [DEBIT:0] score_0_x290;
wire signed [DEBIT:0] score_0_x291;
wire signed [DEBIT:0] score_0_x292;
wire signed [DEBIT:0] score_0_x293;
wire signed [DEBIT:0] score_0_x294;
wire signed [DEBIT:0] score_0_x295;
wire signed [DEBIT:0] score_0_x296;
wire signed [DEBIT:0] score_0_x297;
wire signed [DEBIT:0] score_0_x298;
wire signed [DEBIT:0] score_0_x299;
wire signed [DEBIT:0] score_0_x300;
wire signed [DEBIT:0] score_0_x301;
wire signed [DEBIT:0] score_0_x302;
wire signed [DEBIT:0] score_0_x303;
wire signed [DEBIT:0] score_0_x304;
wire signed [DEBIT:0] score_0_x305;
wire signed [DEBIT:0] score_0_x306;
wire signed [DEBIT:0] score_0_x307;
wire signed [DEBIT:0] score_0_x308;
wire signed [DEBIT:0] score_0_x309;
wire signed [DEBIT:0] score_0_x310;
wire signed [DEBIT:0] score_0_x311;
wire signed [DEBIT:0] score_0_x312;
wire signed [DEBIT:0] score_0_x313;
wire signed [DEBIT:0] score_0_x314;
wire signed [DEBIT:0] score_0_x315;
wire signed [DEBIT:0] score_0_x316;
wire signed [DEBIT:0] score_0_x317;
wire signed [DEBIT:0] score_0_x318;
wire signed [DEBIT:0] score_0_x319;
wire signed [DEBIT:0] score_0_x320;
wire signed [DEBIT:0] score_0_x321;
wire signed [DEBIT:0] score_0_x322;
wire signed [DEBIT:0] score_0_x323;
wire signed [DEBIT:0] score_0_x324;
wire signed [DEBIT:0] score_0_x325;
wire signed [DEBIT:0] score_0_x326;
wire signed [DEBIT:0] score_0_x327;
wire signed [DEBIT:0] score_0_x328;
wire signed [DEBIT:0] score_0_x329;
wire signed [DEBIT:0] score_0_x330;
wire signed [DEBIT:0] score_0_x331;
wire signed [DEBIT:0] score_0_x332;
wire signed [DEBIT:0] score_0_x333;
wire signed [DEBIT:0] score_0_x334;
wire signed [DEBIT:0] score_0_x335;
wire signed [DEBIT:0] score_0_x336;
wire signed [DEBIT:0] score_0_x337;
wire signed [DEBIT:0] score_0_x338;
wire signed [DEBIT:0] score_0_x339;
wire signed [DEBIT:0] score_0_x340;
wire signed [DEBIT:0] score_0_x341;
wire signed [DEBIT:0] score_0_x342;
wire signed [DEBIT:0] score_0_x343;
wire signed [DEBIT:0] score_0_x344;
wire signed [DEBIT:0] score_0_x345;
wire signed [DEBIT:0] score_0_x346;
wire signed [DEBIT:0] score_0_x347;
wire signed [DEBIT:0] score_0_x348;
wire signed [DEBIT:0] score_0_x349;
wire signed [DEBIT:0] score_0_x350;
wire signed [DEBIT:0] score_0_x351;
wire signed [DEBIT:0] score_0_x352;
wire signed [DEBIT:0] score_0_x353;
wire signed [DEBIT:0] score_0_x354;
wire signed [DEBIT:0] score_0_x355;
wire signed [DEBIT:0] score_0_x356;
wire signed [DEBIT:0] score_0_x357;
wire signed [DEBIT:0] score_0_x358;
wire signed [DEBIT:0] score_0_x359;
wire signed [DEBIT:0] score_0_x360;
wire signed [DEBIT:0] score_0_x361;
wire signed [DEBIT:0] score_0_x362;
wire signed [DEBIT:0] score_0_x363;
wire signed [DEBIT:0] score_0_x364;
wire signed [DEBIT:0] score_0_x365;
wire signed [DEBIT:0] score_0_x366;
wire signed [DEBIT:0] score_0_x367;
wire signed [DEBIT:0] score_0_x368;
wire signed [DEBIT:0] score_0_x369;
wire signed [DEBIT:0] score_0_x370;
wire signed [DEBIT:0] score_0_x371;
wire signed [DEBIT:0] score_0_x372;
wire signed [DEBIT:0] score_0_x373;
wire signed [DEBIT:0] score_0_x374;
wire signed [DEBIT:0] score_0_x375;
wire signed [DEBIT:0] score_0_x376;
wire signed [DEBIT:0] score_0_x377;
wire signed [DEBIT:0] score_0_x378;
wire signed [DEBIT:0] score_0_x379;
wire signed [DEBIT:0] score_0_x380;
wire signed [DEBIT:0] score_0_x381;
wire signed [DEBIT:0] score_0_x382;
wire signed [DEBIT:0] score_0_x383;
wire signed [DEBIT:0] score_0_x384;
wire signed [DEBIT:0] score_0_x385;
wire signed [DEBIT:0] score_0_x386;
wire signed [DEBIT:0] score_0_x387;
wire signed [DEBIT:0] score_0_x388;
wire signed [DEBIT:0] score_0_x389;
wire signed [DEBIT:0] score_0_x390;
wire signed [DEBIT:0] score_0_x391;
wire signed [DEBIT:0] score_0_x392;
wire signed [DEBIT:0] score_0_x393;
wire signed [DEBIT:0] score_0_x394;
wire signed [DEBIT:0] score_0_x395;
wire signed [DEBIT:0] score_0_x396;
wire signed [DEBIT:0] score_0_x397;
wire signed [DEBIT:0] score_0_x398;
wire signed [DEBIT:0] score_0_x399;
wire signed [DEBIT:0] score_0_x400;
wire signed [DEBIT:0] score_0_x401;
wire signed [DEBIT:0] score_0_x402;
wire signed [DEBIT:0] score_0_x403;
wire signed [DEBIT:0] score_0_x404;
wire signed [DEBIT:0] score_0_x405;
wire signed [DEBIT:0] score_0_x406;
wire signed [DEBIT:0] score_0_x407;
wire signed [DEBIT:0] score_0_x408;
wire signed [DEBIT:0] score_0_x409;
wire signed [DEBIT:0] score_0_x410;
wire signed [DEBIT:0] score_0_x411;
wire signed [DEBIT:0] score_0_x412;
wire signed [DEBIT:0] score_0_x413;
wire signed [DEBIT:0] score_0_x414;
wire signed [DEBIT:0] score_0_x415;
wire signed [DEBIT:0] score_0_x416;
wire signed [DEBIT:0] score_0_x417;
wire signed [DEBIT:0] score_0_x418;
wire signed [DEBIT:0] score_0_x419;
wire signed [DEBIT:0] score_0_x420;
wire signed [DEBIT:0] score_0_x421;
wire signed [DEBIT:0] score_0_x422;
wire signed [DEBIT:0] score_0_x423;
wire signed [DEBIT:0] score_0_x424;
wire signed [DEBIT:0] score_0_x425;
wire signed [DEBIT:0] score_0_x426;
wire signed [DEBIT:0] score_0_x427;
wire signed [DEBIT:0] score_0_x428;
wire signed [DEBIT:0] score_0_x429;
wire signed [DEBIT:0] score_0_x430;
wire signed [DEBIT:0] score_0_x431;
wire signed [DEBIT:0] score_0_x432;
wire signed [DEBIT:0] score_0_x433;
wire signed [DEBIT:0] score_0_x434;
wire signed [DEBIT:0] score_0_x435;
wire signed [DEBIT:0] score_0_x436;
wire signed [DEBIT:0] score_0_x437;
wire signed [DEBIT:0] score_0_x438;
wire signed [DEBIT:0] score_0_x439;
wire signed [DEBIT:0] score_0_x440;
wire signed [DEBIT:0] score_0_x441;
wire signed [DEBIT:0] score_0_x442;
wire signed [DEBIT:0] score_0_x443;
wire signed [DEBIT:0] score_0_x444;
wire signed [DEBIT:0] score_0_x445;
wire signed [DEBIT:0] score_0_x446;
wire signed [DEBIT:0] score_0_x447;
wire signed [DEBIT:0] score_0_x448;
wire signed [DEBIT:0] score_0_x449;
wire signed [DEBIT:0] score_0_x450;
wire signed [DEBIT:0] score_0_x451;
wire signed [DEBIT:0] score_0_x452;
wire signed [DEBIT:0] score_0_x453;
wire signed [DEBIT:0] score_0_x454;
wire signed [DEBIT:0] score_0_x455;
wire signed [DEBIT:0] score_0_x456;
wire signed [DEBIT:0] score_0_x457;
wire signed [DEBIT:0] score_0_x458;
wire signed [DEBIT:0] score_0_x459;
wire signed [DEBIT:0] score_0_x460;
wire signed [DEBIT:0] score_0_x461;
wire signed [DEBIT:0] score_0_x462;
wire signed [DEBIT:0] score_0_x463;
wire signed [DEBIT:0] score_0_x464;
wire signed [DEBIT:0] score_0_x465;
wire signed [DEBIT:0] score_0_x466;
wire signed [DEBIT:0] score_0_x467;
wire signed [DEBIT:0] score_0_x468;
wire signed [DEBIT:0] score_0_x469;
wire signed [DEBIT:0] score_0_x470;
wire signed [DEBIT:0] score_0_x471;
wire signed [DEBIT:0] score_0_x472;
wire signed [DEBIT:0] score_0_x473;
wire signed [DEBIT:0] score_0_x474;
wire signed [DEBIT:0] score_0_x475;
wire signed [DEBIT:0] score_0_x476;
wire signed [DEBIT:0] score_0_x477;
wire signed [DEBIT:0] score_0_x478;
wire signed [DEBIT:0] score_0_x479;
wire signed [DEBIT:0] score_0_x480;
wire signed [DEBIT:0] score_0_x481;
wire signed [DEBIT:0] score_0_x482;
wire signed [DEBIT:0] score_0_x483;
wire signed [DEBIT:0] score_0_x484;
wire signed [DEBIT:0] score_0_x485;
wire signed [DEBIT:0] score_0_x486;
wire signed [DEBIT:0] score_0_x487;
wire signed [DEBIT:0] score_0_x488;
wire signed [DEBIT:0] score_0_x489;
wire signed [DEBIT:0] score_0_x490;
wire signed [DEBIT:0] score_0_x491;
wire signed [DEBIT:0] score_0_x492;
wire signed [DEBIT:0] score_0_x493;
wire signed [DEBIT:0] score_0_x494;
wire signed [DEBIT:0] score_0_x495;
wire signed [DEBIT:0] score_0_x496;
wire signed [DEBIT:0] score_0_x497;
wire signed [DEBIT:0] score_0_x498;
wire signed [DEBIT:0] score_0_x499;
wire signed [DEBIT:0] score_0_x500;
wire signed [DEBIT:0] score_0_x501;
wire signed [DEBIT:0] score_0_x502;
wire signed [DEBIT:0] score_0_x503;
wire signed [DEBIT:0] score_0_x504;
wire signed [DEBIT:0] score_0_x505;
wire signed [DEBIT:0] score_0_x506;
wire signed [DEBIT:0] score_0_x507;
wire signed [DEBIT:0] score_0_x508;
wire signed [DEBIT:0] score_0_x509;
wire signed [DEBIT:0] score_0_x510;
wire signed [DEBIT:0] score_0_x511;
wire signed [DEBIT:0] score_0_x512;
wire signed [DEBIT:0] score_0_x513;
wire signed [DEBIT:0] score_0_x514;
wire signed [DEBIT:0] score_0_x515;
wire signed [DEBIT:0] score_0_x516;
wire signed [DEBIT:0] score_0_x517;
wire signed [DEBIT:0] score_0_x518;
wire signed [DEBIT:0] score_0_x519;
wire signed [DEBIT:0] score_0_x520;
wire signed [DEBIT:0] score_0_x521;
wire signed [DEBIT:0] score_0_x522;
wire signed [DEBIT:0] score_0_x523;
wire signed [DEBIT:0] score_0_x524;
wire signed [DEBIT:0] score_0_x525;
wire signed [DEBIT:0] score_0_x526;
wire signed [DEBIT:0] score_0_x527;
wire signed [DEBIT:0] score_0_x528;
wire signed [DEBIT:0] score_0_x529;
wire signed [DEBIT:0] score_0_x530;
wire signed [DEBIT:0] score_0_x531;
wire signed [DEBIT:0] score_0_x532;
wire signed [DEBIT:0] score_0_x533;
wire signed [DEBIT:0] score_0_x534;
wire signed [DEBIT:0] score_0_x535;
wire signed [DEBIT:0] score_0_x536;
wire signed [DEBIT:0] score_0_x537;
wire signed [DEBIT:0] score_0_x538;
wire signed [DEBIT:0] score_0_x539;
wire signed [DEBIT:0] score_0_x540;
wire signed [DEBIT:0] score_0_x541;
wire signed [DEBIT:0] score_0_x542;
wire signed [DEBIT:0] score_0_x543;
wire signed [DEBIT:0] score_0_x544;
wire signed [DEBIT:0] score_0_x545;
wire signed [DEBIT:0] score_0_x546;
wire signed [DEBIT:0] score_0_x547;
wire signed [DEBIT:0] score_0_x548;
wire signed [DEBIT:0] score_0_x549;
wire signed [DEBIT:0] score_0_x550;
wire signed [DEBIT:0] score_0_x551;
wire signed [DEBIT:0] score_0_x552;
wire signed [DEBIT:0] score_0_x553;
wire signed [DEBIT:0] score_0_x554;
wire signed [DEBIT:0] score_0_x555;
wire signed [DEBIT:0] score_0_x556;
wire signed [DEBIT:0] score_0_x557;
wire signed [DEBIT:0] score_0_x558;
wire signed [DEBIT:0] score_0_x559;
wire signed [DEBIT:0] score_0_x560;
wire signed [DEBIT:0] score_0_x561;
wire signed [DEBIT:0] score_0_x562;
wire signed [DEBIT:0] score_0_x563;
wire signed [DEBIT:0] score_0_x564;
wire signed [DEBIT:0] score_0_x565;
wire signed [DEBIT:0] score_0_x566;
wire signed [DEBIT:0] score_0_x567;
wire signed [DEBIT:0] score_0_x568;
wire signed [DEBIT:0] score_0_x569;
wire signed [DEBIT:0] score_0_x570;
wire signed [DEBIT:0] score_0_x571;
wire signed [DEBIT:0] score_0_x572;
wire signed [DEBIT:0] score_0_x573;
wire signed [DEBIT:0] score_0_x574;
wire signed [DEBIT:0] score_0_x575;
wire signed [DEBIT:0] score_0_x576;
wire signed [DEBIT:0] score_0_x577;
wire signed [DEBIT:0] score_0_x578;
wire signed [DEBIT:0] score_0_x579;
wire signed [DEBIT:0] score_0_x580;
wire signed [DEBIT:0] score_0_x581;
wire signed [DEBIT:0] score_0_x582;
wire signed [DEBIT:0] score_0_x583;
wire signed [DEBIT:0] score_0_x584;
wire signed [DEBIT:0] score_0_x585;
wire signed [DEBIT:0] score_0_x586;
wire signed [DEBIT:0] score_0_x587;
wire signed [DEBIT:0] score_0_x588;
wire signed [DEBIT:0] score_0_x589;
wire signed [DEBIT:0] score_0_x590;
wire signed [DEBIT:0] score_0_x591;
wire signed [DEBIT:0] score_0_x592;
wire signed [DEBIT:0] score_0_x593;
wire signed [DEBIT:0] score_0_x594;
wire signed [DEBIT:0] score_0_x595;
wire signed [DEBIT:0] score_0_x596;
wire signed [DEBIT:0] score_0_x597;
wire signed [DEBIT:0] score_0_x598;
wire signed [DEBIT:0] score_0_x599;
wire signed [DEBIT:0] score_0_x600;
wire signed [DEBIT:0] score_0_x601;
wire signed [DEBIT:0] score_0_x602;
wire signed [DEBIT:0] score_0_x603;
wire signed [DEBIT:0] score_0_x604;
wire signed [DEBIT:0] score_0_x605;
wire signed [DEBIT:0] score_0_x606;
wire signed [DEBIT:0] score_0_x607;
wire signed [DEBIT:0] score_0_x608;
wire signed [DEBIT:0] score_0_x609;
wire signed [DEBIT:0] score_0_x610;
wire signed [DEBIT:0] score_0_x611;
wire signed [DEBIT:0] score_0_x612;
wire signed [DEBIT:0] score_0_x613;
wire signed [DEBIT:0] score_0_x614;
wire signed [DEBIT:0] score_0_x615;
wire signed [DEBIT:0] score_0_x616;
wire signed [DEBIT:0] score_0_x617;
wire signed [DEBIT:0] score_0_x618;
wire signed [DEBIT:0] score_0_x619;
wire signed [DEBIT:0] score_0_x620;
wire signed [DEBIT:0] score_0_x621;
wire signed [DEBIT:0] score_0_x622;
wire signed [DEBIT:0] score_0_x623;
wire signed [DEBIT:0] score_0_x624;
wire signed [DEBIT:0] score_0_x625;
wire signed [DEBIT:0] score_0_x626;
wire signed [DEBIT:0] score_0_x627;
wire signed [DEBIT:0] score_0_x628;
wire signed [DEBIT:0] score_0_x629;
wire signed [DEBIT:0] score_0_x630;
wire signed [DEBIT:0] score_0_x631;
wire signed [DEBIT:0] score_0_x632;
wire signed [DEBIT:0] score_0_x633;
wire signed [DEBIT:0] score_0_x634;
wire signed [DEBIT:0] score_0_x635;
wire signed [DEBIT:0] score_0_x636;
wire signed [DEBIT:0] score_0_x637;
wire signed [DEBIT:0] score_0_x638;
wire signed [DEBIT:0] score_0_x639;
wire signed [DEBIT:0] score_0_x640;
wire signed [DEBIT:0] score_0_x641;
wire signed [DEBIT:0] score_0_x642;
wire signed [DEBIT:0] score_0_x643;
wire signed [DEBIT:0] score_0_x644;
wire signed [DEBIT:0] score_0_x645;
wire signed [DEBIT:0] score_0_x646;
wire signed [DEBIT:0] score_0_x647;
wire signed [DEBIT:0] score_0_x648;
wire signed [DEBIT:0] score_0_x649;
wire signed [DEBIT:0] score_0_x650;
wire signed [DEBIT:0] score_0_x651;
wire signed [DEBIT:0] score_0_x652;
wire signed [DEBIT:0] score_0_x653;
wire signed [DEBIT:0] score_0_x654;
wire signed [DEBIT:0] score_0_x655;
wire signed [DEBIT:0] score_0_x656;
wire signed [DEBIT:0] score_0_x657;
wire signed [DEBIT:0] score_0_x658;
wire signed [DEBIT:0] score_0_x659;
wire signed [DEBIT:0] score_0_x660;
wire signed [DEBIT:0] score_0_x661;
wire signed [DEBIT:0] score_0_x662;
wire signed [DEBIT:0] score_0_x663;
wire signed [DEBIT:0] score_0_x664;
wire signed [DEBIT:0] score_0_x665;
wire signed [DEBIT:0] score_0_x666;
wire signed [DEBIT:0] score_0_x667;
wire signed [DEBIT:0] score_0_x668;
wire signed [DEBIT:0] score_0_x669;
wire signed [DEBIT:0] score_0_x670;
wire signed [DEBIT:0] score_0_x671;
wire signed [DEBIT:0] score_0_x672;
wire signed [DEBIT:0] score_0_x673;
wire signed [DEBIT:0] score_0_x674;
wire signed [DEBIT:0] score_0_x675;
wire signed [DEBIT:0] score_0_x676;
wire signed [DEBIT:0] score_0_x677;
wire signed [DEBIT:0] score_0_x678;
wire signed [DEBIT:0] score_0_x679;
wire signed [DEBIT:0] score_0_x680;
wire signed [DEBIT:0] score_0_x681;
wire signed [DEBIT:0] score_0_x682;
wire signed [DEBIT:0] score_0_x683;
wire signed [DEBIT:0] score_0_x684;
wire signed [DEBIT:0] score_0_x685;
wire signed [DEBIT:0] score_0_x686;
wire signed [DEBIT:0] score_0_x687;
wire signed [DEBIT:0] score_0_x688;
wire signed [DEBIT:0] score_0_x689;
wire signed [DEBIT:0] score_0_x690;
wire signed [DEBIT:0] score_0_x691;
wire signed [DEBIT:0] score_0_x692;
wire signed [DEBIT:0] score_0_x693;
wire signed [DEBIT:0] score_0_x694;
wire signed [DEBIT:0] score_0_x695;
wire signed [DEBIT:0] score_0_x696;
wire signed [DEBIT:0] score_0_x697;
wire signed [DEBIT:0] score_0_x698;
wire signed [DEBIT:0] score_0_x699;
wire signed [DEBIT:0] score_0_x700;
wire signed [DEBIT:0] score_0_x701;
wire signed [DEBIT:0] score_0_x702;
wire signed [DEBIT:0] score_0_x703;
wire signed [DEBIT:0] score_0_x704;
wire signed [DEBIT:0] score_0_x705;
wire signed [DEBIT:0] score_0_x706;
wire signed [DEBIT:0] score_0_x707;
wire signed [DEBIT:0] score_0_x708;
wire signed [DEBIT:0] score_0_x709;
wire signed [DEBIT:0] score_0_x710;
wire signed [DEBIT:0] score_0_x711;
wire signed [DEBIT:0] score_0_x712;
wire signed [DEBIT:0] score_0_x713;
wire signed [DEBIT:0] score_0_x714;
wire signed [DEBIT:0] score_0_x715;
wire signed [DEBIT:0] score_0_x716;
wire signed [DEBIT:0] score_0_x717;
wire signed [DEBIT:0] score_0_x718;
wire signed [DEBIT:0] score_0_x719;
wire signed [DEBIT:0] score_0_x720;
wire signed [DEBIT:0] score_0_x721;
wire signed [DEBIT:0] score_0_x722;
wire signed [DEBIT:0] score_0_x723;
wire signed [DEBIT:0] score_0_x724;
wire signed [DEBIT:0] score_0_x725;
wire signed [DEBIT:0] score_0_x726;
wire signed [DEBIT:0] score_0_x727;
wire signed [DEBIT:0] score_0_x728;
wire signed [DEBIT:0] score_0_x729;
wire signed [DEBIT:0] score_0_x730;
wire signed [DEBIT:0] score_0_x731;
wire signed [DEBIT:0] score_0_x732;
wire signed [DEBIT:0] score_0_x733;
wire signed [DEBIT:0] score_0_x734;
wire signed [DEBIT:0] score_0_x735;
wire signed [DEBIT:0] score_0_x736;
wire signed [DEBIT:0] score_0_x737;
wire signed [DEBIT:0] score_0_x738;
wire signed [DEBIT:0] score_0_x739;
wire signed [DEBIT:0] score_0_x740;
wire signed [DEBIT:0] score_0_x741;
wire signed [DEBIT:0] score_0_x742;
wire signed [DEBIT:0] score_0_x743;
wire signed [DEBIT:0] score_0_x744;
wire signed [DEBIT:0] score_0_x745;
wire signed [DEBIT:0] score_0_x746;
wire signed [DEBIT:0] score_0_x747;
wire signed [DEBIT:0] score_0_x748;
wire signed [DEBIT:0] score_0_x749;
wire signed [DEBIT:0] score_0_x750;
wire signed [DEBIT:0] score_0_x751;
wire signed [DEBIT:0] score_0_x752;
wire signed [DEBIT:0] score_0_x753;
wire signed [DEBIT:0] score_0_x754;
wire signed [DEBIT:0] score_0_x755;
wire signed [DEBIT:0] score_0_x756;
wire signed [DEBIT:0] score_0_x757;
wire signed [DEBIT:0] score_0_x758;
wire signed [DEBIT:0] score_0_x759;
wire signed [DEBIT:0] score_0_x760;
wire signed [DEBIT:0] score_0_x761;
wire signed [DEBIT:0] score_0_x762;
wire signed [DEBIT:0] score_0_x763;
wire signed [DEBIT:0] score_0_x764;
wire signed [DEBIT:0] score_0_x765;
wire signed [DEBIT:0] score_0_x766;
wire signed [DEBIT:0] score_0_x767;
wire signed [DEBIT:0] score_0_x768;
wire signed [DEBIT:0] score_0_x769;
wire signed [DEBIT:0] score_0_x770;
wire signed [DEBIT:0] score_0_x771;
wire signed [DEBIT:0] score_0_x772;
wire signed [DEBIT:0] score_0_x773;
wire signed [DEBIT:0] score_0_x774;
wire signed [DEBIT:0] score_0_x775;
wire signed [DEBIT:0] score_0_x776;
wire signed [DEBIT:0] score_0_x777;
wire signed [DEBIT:0] score_0_x778;
wire signed [DEBIT:0] score_0_x779;
wire signed [DEBIT:0] score_0_x780;
wire signed [DEBIT:0] score_0_x781;
wire signed [DEBIT:0] score_0_x782;
wire signed [DEBIT:0] score_0_x783;
wire signed [DEBIT:0] score_0_x784;
wire signed [DEBIT:0] score_1_x1;
wire signed [DEBIT:0] score_1_x2;
wire signed [DEBIT:0] score_1_x3;
wire signed [DEBIT:0] score_1_x4;
wire signed [DEBIT:0] score_1_x5;
wire signed [DEBIT:0] score_1_x6;
wire signed [DEBIT:0] score_1_x7;
wire signed [DEBIT:0] score_1_x8;
wire signed [DEBIT:0] score_1_x9;
wire signed [DEBIT:0] score_1_x10;
wire signed [DEBIT:0] score_1_x11;
wire signed [DEBIT:0] score_1_x12;
wire signed [DEBIT:0] score_1_x13;
wire signed [DEBIT:0] score_1_x14;
wire signed [DEBIT:0] score_1_x15;
wire signed [DEBIT:0] score_1_x16;
wire signed [DEBIT:0] score_1_x17;
wire signed [DEBIT:0] score_1_x18;
wire signed [DEBIT:0] score_1_x19;
wire signed [DEBIT:0] score_1_x20;
wire signed [DEBIT:0] score_1_x21;
wire signed [DEBIT:0] score_1_x22;
wire signed [DEBIT:0] score_1_x23;
wire signed [DEBIT:0] score_1_x24;
wire signed [DEBIT:0] score_1_x25;
wire signed [DEBIT:0] score_1_x26;
wire signed [DEBIT:0] score_1_x27;
wire signed [DEBIT:0] score_1_x28;
wire signed [DEBIT:0] score_1_x29;
wire signed [DEBIT:0] score_1_x30;
wire signed [DEBIT:0] score_1_x31;
wire signed [DEBIT:0] score_1_x32;
wire signed [DEBIT:0] score_1_x33;
wire signed [DEBIT:0] score_1_x34;
wire signed [DEBIT:0] score_1_x35;
wire signed [DEBIT:0] score_1_x36;
wire signed [DEBIT:0] score_1_x37;
wire signed [DEBIT:0] score_1_x38;
wire signed [DEBIT:0] score_1_x39;
wire signed [DEBIT:0] score_1_x40;
wire signed [DEBIT:0] score_1_x41;
wire signed [DEBIT:0] score_1_x42;
wire signed [DEBIT:0] score_1_x43;
wire signed [DEBIT:0] score_1_x44;
wire signed [DEBIT:0] score_1_x45;
wire signed [DEBIT:0] score_1_x46;
wire signed [DEBIT:0] score_1_x47;
wire signed [DEBIT:0] score_1_x48;
wire signed [DEBIT:0] score_1_x49;
wire signed [DEBIT:0] score_1_x50;
wire signed [DEBIT:0] score_1_x51;
wire signed [DEBIT:0] score_1_x52;
wire signed [DEBIT:0] score_1_x53;
wire signed [DEBIT:0] score_1_x54;
wire signed [DEBIT:0] score_1_x55;
wire signed [DEBIT:0] score_1_x56;
wire signed [DEBIT:0] score_1_x57;
wire signed [DEBIT:0] score_1_x58;
wire signed [DEBIT:0] score_1_x59;
wire signed [DEBIT:0] score_1_x60;
wire signed [DEBIT:0] score_1_x61;
wire signed [DEBIT:0] score_1_x62;
wire signed [DEBIT:0] score_1_x63;
wire signed [DEBIT:0] score_1_x64;
wire signed [DEBIT:0] score_1_x65;
wire signed [DEBIT:0] score_1_x66;
wire signed [DEBIT:0] score_1_x67;
wire signed [DEBIT:0] score_1_x68;
wire signed [DEBIT:0] score_1_x69;
wire signed [DEBIT:0] score_1_x70;
wire signed [DEBIT:0] score_1_x71;
wire signed [DEBIT:0] score_1_x72;
wire signed [DEBIT:0] score_1_x73;
wire signed [DEBIT:0] score_1_x74;
wire signed [DEBIT:0] score_1_x75;
wire signed [DEBIT:0] score_1_x76;
wire signed [DEBIT:0] score_1_x77;
wire signed [DEBIT:0] score_1_x78;
wire signed [DEBIT:0] score_1_x79;
wire signed [DEBIT:0] score_1_x80;
wire signed [DEBIT:0] score_1_x81;
wire signed [DEBIT:0] score_1_x82;
wire signed [DEBIT:0] score_1_x83;
wire signed [DEBIT:0] score_1_x84;
wire signed [DEBIT:0] score_1_x85;
wire signed [DEBIT:0] score_1_x86;
wire signed [DEBIT:0] score_1_x87;
wire signed [DEBIT:0] score_1_x88;
wire signed [DEBIT:0] score_1_x89;
wire signed [DEBIT:0] score_1_x90;
wire signed [DEBIT:0] score_1_x91;
wire signed [DEBIT:0] score_1_x92;
wire signed [DEBIT:0] score_1_x93;
wire signed [DEBIT:0] score_1_x94;
wire signed [DEBIT:0] score_1_x95;
wire signed [DEBIT:0] score_1_x96;
wire signed [DEBIT:0] score_1_x97;
wire signed [DEBIT:0] score_1_x98;
wire signed [DEBIT:0] score_1_x99;
wire signed [DEBIT:0] score_1_x100;
wire signed [DEBIT:0] score_1_x101;
wire signed [DEBIT:0] score_1_x102;
wire signed [DEBIT:0] score_1_x103;
wire signed [DEBIT:0] score_1_x104;
wire signed [DEBIT:0] score_1_x105;
wire signed [DEBIT:0] score_1_x106;
wire signed [DEBIT:0] score_1_x107;
wire signed [DEBIT:0] score_1_x108;
wire signed [DEBIT:0] score_1_x109;
wire signed [DEBIT:0] score_1_x110;
wire signed [DEBIT:0] score_1_x111;
wire signed [DEBIT:0] score_1_x112;
wire signed [DEBIT:0] score_1_x113;
wire signed [DEBIT:0] score_1_x114;
wire signed [DEBIT:0] score_1_x115;
wire signed [DEBIT:0] score_1_x116;
wire signed [DEBIT:0] score_1_x117;
wire signed [DEBIT:0] score_1_x118;
wire signed [DEBIT:0] score_1_x119;
wire signed [DEBIT:0] score_1_x120;
wire signed [DEBIT:0] score_1_x121;
wire signed [DEBIT:0] score_1_x122;
wire signed [DEBIT:0] score_1_x123;
wire signed [DEBIT:0] score_1_x124;
wire signed [DEBIT:0] score_1_x125;
wire signed [DEBIT:0] score_1_x126;
wire signed [DEBIT:0] score_1_x127;
wire signed [DEBIT:0] score_1_x128;
wire signed [DEBIT:0] score_1_x129;
wire signed [DEBIT:0] score_1_x130;
wire signed [DEBIT:0] score_1_x131;
wire signed [DEBIT:0] score_1_x132;
wire signed [DEBIT:0] score_1_x133;
wire signed [DEBIT:0] score_1_x134;
wire signed [DEBIT:0] score_1_x135;
wire signed [DEBIT:0] score_1_x136;
wire signed [DEBIT:0] score_1_x137;
wire signed [DEBIT:0] score_1_x138;
wire signed [DEBIT:0] score_1_x139;
wire signed [DEBIT:0] score_1_x140;
wire signed [DEBIT:0] score_1_x141;
wire signed [DEBIT:0] score_1_x142;
wire signed [DEBIT:0] score_1_x143;
wire signed [DEBIT:0] score_1_x144;
wire signed [DEBIT:0] score_1_x145;
wire signed [DEBIT:0] score_1_x146;
wire signed [DEBIT:0] score_1_x147;
wire signed [DEBIT:0] score_1_x148;
wire signed [DEBIT:0] score_1_x149;
wire signed [DEBIT:0] score_1_x150;
wire signed [DEBIT:0] score_1_x151;
wire signed [DEBIT:0] score_1_x152;
wire signed [DEBIT:0] score_1_x153;
wire signed [DEBIT:0] score_1_x154;
wire signed [DEBIT:0] score_1_x155;
wire signed [DEBIT:0] score_1_x156;
wire signed [DEBIT:0] score_1_x157;
wire signed [DEBIT:0] score_1_x158;
wire signed [DEBIT:0] score_1_x159;
wire signed [DEBIT:0] score_1_x160;
wire signed [DEBIT:0] score_1_x161;
wire signed [DEBIT:0] score_1_x162;
wire signed [DEBIT:0] score_1_x163;
wire signed [DEBIT:0] score_1_x164;
wire signed [DEBIT:0] score_1_x165;
wire signed [DEBIT:0] score_1_x166;
wire signed [DEBIT:0] score_1_x167;
wire signed [DEBIT:0] score_1_x168;
wire signed [DEBIT:0] score_1_x169;
wire signed [DEBIT:0] score_1_x170;
wire signed [DEBIT:0] score_1_x171;
wire signed [DEBIT:0] score_1_x172;
wire signed [DEBIT:0] score_1_x173;
wire signed [DEBIT:0] score_1_x174;
wire signed [DEBIT:0] score_1_x175;
wire signed [DEBIT:0] score_1_x176;
wire signed [DEBIT:0] score_1_x177;
wire signed [DEBIT:0] score_1_x178;
wire signed [DEBIT:0] score_1_x179;
wire signed [DEBIT:0] score_1_x180;
wire signed [DEBIT:0] score_1_x181;
wire signed [DEBIT:0] score_1_x182;
wire signed [DEBIT:0] score_1_x183;
wire signed [DEBIT:0] score_1_x184;
wire signed [DEBIT:0] score_1_x185;
wire signed [DEBIT:0] score_1_x186;
wire signed [DEBIT:0] score_1_x187;
wire signed [DEBIT:0] score_1_x188;
wire signed [DEBIT:0] score_1_x189;
wire signed [DEBIT:0] score_1_x190;
wire signed [DEBIT:0] score_1_x191;
wire signed [DEBIT:0] score_1_x192;
wire signed [DEBIT:0] score_1_x193;
wire signed [DEBIT:0] score_1_x194;
wire signed [DEBIT:0] score_1_x195;
wire signed [DEBIT:0] score_1_x196;
wire signed [DEBIT:0] score_1_x197;
wire signed [DEBIT:0] score_1_x198;
wire signed [DEBIT:0] score_1_x199;
wire signed [DEBIT:0] score_1_x200;
wire signed [DEBIT:0] score_1_x201;
wire signed [DEBIT:0] score_1_x202;
wire signed [DEBIT:0] score_1_x203;
wire signed [DEBIT:0] score_1_x204;
wire signed [DEBIT:0] score_1_x205;
wire signed [DEBIT:0] score_1_x206;
wire signed [DEBIT:0] score_1_x207;
wire signed [DEBIT:0] score_1_x208;
wire signed [DEBIT:0] score_1_x209;
wire signed [DEBIT:0] score_1_x210;
wire signed [DEBIT:0] score_1_x211;
wire signed [DEBIT:0] score_1_x212;
wire signed [DEBIT:0] score_1_x213;
wire signed [DEBIT:0] score_1_x214;
wire signed [DEBIT:0] score_1_x215;
wire signed [DEBIT:0] score_1_x216;
wire signed [DEBIT:0] score_1_x217;
wire signed [DEBIT:0] score_1_x218;
wire signed [DEBIT:0] score_1_x219;
wire signed [DEBIT:0] score_1_x220;
wire signed [DEBIT:0] score_1_x221;
wire signed [DEBIT:0] score_1_x222;
wire signed [DEBIT:0] score_1_x223;
wire signed [DEBIT:0] score_1_x224;
wire signed [DEBIT:0] score_1_x225;
wire signed [DEBIT:0] score_1_x226;
wire signed [DEBIT:0] score_1_x227;
wire signed [DEBIT:0] score_1_x228;
wire signed [DEBIT:0] score_1_x229;
wire signed [DEBIT:0] score_1_x230;
wire signed [DEBIT:0] score_1_x231;
wire signed [DEBIT:0] score_1_x232;
wire signed [DEBIT:0] score_1_x233;
wire signed [DEBIT:0] score_1_x234;
wire signed [DEBIT:0] score_1_x235;
wire signed [DEBIT:0] score_1_x236;
wire signed [DEBIT:0] score_1_x237;
wire signed [DEBIT:0] score_1_x238;
wire signed [DEBIT:0] score_1_x239;
wire signed [DEBIT:0] score_1_x240;
wire signed [DEBIT:0] score_1_x241;
wire signed [DEBIT:0] score_1_x242;
wire signed [DEBIT:0] score_1_x243;
wire signed [DEBIT:0] score_1_x244;
wire signed [DEBIT:0] score_1_x245;
wire signed [DEBIT:0] score_1_x246;
wire signed [DEBIT:0] score_1_x247;
wire signed [DEBIT:0] score_1_x248;
wire signed [DEBIT:0] score_1_x249;
wire signed [DEBIT:0] score_1_x250;
wire signed [DEBIT:0] score_1_x251;
wire signed [DEBIT:0] score_1_x252;
wire signed [DEBIT:0] score_1_x253;
wire signed [DEBIT:0] score_1_x254;
wire signed [DEBIT:0] score_1_x255;
wire signed [DEBIT:0] score_1_x256;
wire signed [DEBIT:0] score_1_x257;
wire signed [DEBIT:0] score_1_x258;
wire signed [DEBIT:0] score_1_x259;
wire signed [DEBIT:0] score_1_x260;
wire signed [DEBIT:0] score_1_x261;
wire signed [DEBIT:0] score_1_x262;
wire signed [DEBIT:0] score_1_x263;
wire signed [DEBIT:0] score_1_x264;
wire signed [DEBIT:0] score_1_x265;
wire signed [DEBIT:0] score_1_x266;
wire signed [DEBIT:0] score_1_x267;
wire signed [DEBIT:0] score_1_x268;
wire signed [DEBIT:0] score_1_x269;
wire signed [DEBIT:0] score_1_x270;
wire signed [DEBIT:0] score_1_x271;
wire signed [DEBIT:0] score_1_x272;
wire signed [DEBIT:0] score_1_x273;
wire signed [DEBIT:0] score_1_x274;
wire signed [DEBIT:0] score_1_x275;
wire signed [DEBIT:0] score_1_x276;
wire signed [DEBIT:0] score_1_x277;
wire signed [DEBIT:0] score_1_x278;
wire signed [DEBIT:0] score_1_x279;
wire signed [DEBIT:0] score_1_x280;
wire signed [DEBIT:0] score_1_x281;
wire signed [DEBIT:0] score_1_x282;
wire signed [DEBIT:0] score_1_x283;
wire signed [DEBIT:0] score_1_x284;
wire signed [DEBIT:0] score_1_x285;
wire signed [DEBIT:0] score_1_x286;
wire signed [DEBIT:0] score_1_x287;
wire signed [DEBIT:0] score_1_x288;
wire signed [DEBIT:0] score_1_x289;
wire signed [DEBIT:0] score_1_x290;
wire signed [DEBIT:0] score_1_x291;
wire signed [DEBIT:0] score_1_x292;
wire signed [DEBIT:0] score_1_x293;
wire signed [DEBIT:0] score_1_x294;
wire signed [DEBIT:0] score_1_x295;
wire signed [DEBIT:0] score_1_x296;
wire signed [DEBIT:0] score_1_x297;
wire signed [DEBIT:0] score_1_x298;
wire signed [DEBIT:0] score_1_x299;
wire signed [DEBIT:0] score_1_x300;
wire signed [DEBIT:0] score_1_x301;
wire signed [DEBIT:0] score_1_x302;
wire signed [DEBIT:0] score_1_x303;
wire signed [DEBIT:0] score_1_x304;
wire signed [DEBIT:0] score_1_x305;
wire signed [DEBIT:0] score_1_x306;
wire signed [DEBIT:0] score_1_x307;
wire signed [DEBIT:0] score_1_x308;
wire signed [DEBIT:0] score_1_x309;
wire signed [DEBIT:0] score_1_x310;
wire signed [DEBIT:0] score_1_x311;
wire signed [DEBIT:0] score_1_x312;
wire signed [DEBIT:0] score_1_x313;
wire signed [DEBIT:0] score_1_x314;
wire signed [DEBIT:0] score_1_x315;
wire signed [DEBIT:0] score_1_x316;
wire signed [DEBIT:0] score_1_x317;
wire signed [DEBIT:0] score_1_x318;
wire signed [DEBIT:0] score_1_x319;
wire signed [DEBIT:0] score_1_x320;
wire signed [DEBIT:0] score_1_x321;
wire signed [DEBIT:0] score_1_x322;
wire signed [DEBIT:0] score_1_x323;
wire signed [DEBIT:0] score_1_x324;
wire signed [DEBIT:0] score_1_x325;
wire signed [DEBIT:0] score_1_x326;
wire signed [DEBIT:0] score_1_x327;
wire signed [DEBIT:0] score_1_x328;
wire signed [DEBIT:0] score_1_x329;
wire signed [DEBIT:0] score_1_x330;
wire signed [DEBIT:0] score_1_x331;
wire signed [DEBIT:0] score_1_x332;
wire signed [DEBIT:0] score_1_x333;
wire signed [DEBIT:0] score_1_x334;
wire signed [DEBIT:0] score_1_x335;
wire signed [DEBIT:0] score_1_x336;
wire signed [DEBIT:0] score_1_x337;
wire signed [DEBIT:0] score_1_x338;
wire signed [DEBIT:0] score_1_x339;
wire signed [DEBIT:0] score_1_x340;
wire signed [DEBIT:0] score_1_x341;
wire signed [DEBIT:0] score_1_x342;
wire signed [DEBIT:0] score_1_x343;
wire signed [DEBIT:0] score_1_x344;
wire signed [DEBIT:0] score_1_x345;
wire signed [DEBIT:0] score_1_x346;
wire signed [DEBIT:0] score_1_x347;
wire signed [DEBIT:0] score_1_x348;
wire signed [DEBIT:0] score_1_x349;
wire signed [DEBIT:0] score_1_x350;
wire signed [DEBIT:0] score_1_x351;
wire signed [DEBIT:0] score_1_x352;
wire signed [DEBIT:0] score_1_x353;
wire signed [DEBIT:0] score_1_x354;
wire signed [DEBIT:0] score_1_x355;
wire signed [DEBIT:0] score_1_x356;
wire signed [DEBIT:0] score_1_x357;
wire signed [DEBIT:0] score_1_x358;
wire signed [DEBIT:0] score_1_x359;
wire signed [DEBIT:0] score_1_x360;
wire signed [DEBIT:0] score_1_x361;
wire signed [DEBIT:0] score_1_x362;
wire signed [DEBIT:0] score_1_x363;
wire signed [DEBIT:0] score_1_x364;
wire signed [DEBIT:0] score_1_x365;
wire signed [DEBIT:0] score_1_x366;
wire signed [DEBIT:0] score_1_x367;
wire signed [DEBIT:0] score_1_x368;
wire signed [DEBIT:0] score_1_x369;
wire signed [DEBIT:0] score_1_x370;
wire signed [DEBIT:0] score_1_x371;
wire signed [DEBIT:0] score_1_x372;
wire signed [DEBIT:0] score_1_x373;
wire signed [DEBIT:0] score_1_x374;
wire signed [DEBIT:0] score_1_x375;
wire signed [DEBIT:0] score_1_x376;
wire signed [DEBIT:0] score_1_x377;
wire signed [DEBIT:0] score_1_x378;
wire signed [DEBIT:0] score_1_x379;
wire signed [DEBIT:0] score_1_x380;
wire signed [DEBIT:0] score_1_x381;
wire signed [DEBIT:0] score_1_x382;
wire signed [DEBIT:0] score_1_x383;
wire signed [DEBIT:0] score_1_x384;
wire signed [DEBIT:0] score_1_x385;
wire signed [DEBIT:0] score_1_x386;
wire signed [DEBIT:0] score_1_x387;
wire signed [DEBIT:0] score_1_x388;
wire signed [DEBIT:0] score_1_x389;
wire signed [DEBIT:0] score_1_x390;
wire signed [DEBIT:0] score_1_x391;
wire signed [DEBIT:0] score_1_x392;
wire signed [DEBIT:0] score_1_x393;
wire signed [DEBIT:0] score_1_x394;
wire signed [DEBIT:0] score_1_x395;
wire signed [DEBIT:0] score_1_x396;
wire signed [DEBIT:0] score_1_x397;
wire signed [DEBIT:0] score_1_x398;
wire signed [DEBIT:0] score_1_x399;
wire signed [DEBIT:0] score_1_x400;
wire signed [DEBIT:0] score_1_x401;
wire signed [DEBIT:0] score_1_x402;
wire signed [DEBIT:0] score_1_x403;
wire signed [DEBIT:0] score_1_x404;
wire signed [DEBIT:0] score_1_x405;
wire signed [DEBIT:0] score_1_x406;
wire signed [DEBIT:0] score_1_x407;
wire signed [DEBIT:0] score_1_x408;
wire signed [DEBIT:0] score_1_x409;
wire signed [DEBIT:0] score_1_x410;
wire signed [DEBIT:0] score_1_x411;
wire signed [DEBIT:0] score_1_x412;
wire signed [DEBIT:0] score_1_x413;
wire signed [DEBIT:0] score_1_x414;
wire signed [DEBIT:0] score_1_x415;
wire signed [DEBIT:0] score_1_x416;
wire signed [DEBIT:0] score_1_x417;
wire signed [DEBIT:0] score_1_x418;
wire signed [DEBIT:0] score_1_x419;
wire signed [DEBIT:0] score_1_x420;
wire signed [DEBIT:0] score_1_x421;
wire signed [DEBIT:0] score_1_x422;
wire signed [DEBIT:0] score_1_x423;
wire signed [DEBIT:0] score_1_x424;
wire signed [DEBIT:0] score_1_x425;
wire signed [DEBIT:0] score_1_x426;
wire signed [DEBIT:0] score_1_x427;
wire signed [DEBIT:0] score_1_x428;
wire signed [DEBIT:0] score_1_x429;
wire signed [DEBIT:0] score_1_x430;
wire signed [DEBIT:0] score_1_x431;
wire signed [DEBIT:0] score_1_x432;
wire signed [DEBIT:0] score_1_x433;
wire signed [DEBIT:0] score_1_x434;
wire signed [DEBIT:0] score_1_x435;
wire signed [DEBIT:0] score_1_x436;
wire signed [DEBIT:0] score_1_x437;
wire signed [DEBIT:0] score_1_x438;
wire signed [DEBIT:0] score_1_x439;
wire signed [DEBIT:0] score_1_x440;
wire signed [DEBIT:0] score_1_x441;
wire signed [DEBIT:0] score_1_x442;
wire signed [DEBIT:0] score_1_x443;
wire signed [DEBIT:0] score_1_x444;
wire signed [DEBIT:0] score_1_x445;
wire signed [DEBIT:0] score_1_x446;
wire signed [DEBIT:0] score_1_x447;
wire signed [DEBIT:0] score_1_x448;
wire signed [DEBIT:0] score_1_x449;
wire signed [DEBIT:0] score_1_x450;
wire signed [DEBIT:0] score_1_x451;
wire signed [DEBIT:0] score_1_x452;
wire signed [DEBIT:0] score_1_x453;
wire signed [DEBIT:0] score_1_x454;
wire signed [DEBIT:0] score_1_x455;
wire signed [DEBIT:0] score_1_x456;
wire signed [DEBIT:0] score_1_x457;
wire signed [DEBIT:0] score_1_x458;
wire signed [DEBIT:0] score_1_x459;
wire signed [DEBIT:0] score_1_x460;
wire signed [DEBIT:0] score_1_x461;
wire signed [DEBIT:0] score_1_x462;
wire signed [DEBIT:0] score_1_x463;
wire signed [DEBIT:0] score_1_x464;
wire signed [DEBIT:0] score_1_x465;
wire signed [DEBIT:0] score_1_x466;
wire signed [DEBIT:0] score_1_x467;
wire signed [DEBIT:0] score_1_x468;
wire signed [DEBIT:0] score_1_x469;
wire signed [DEBIT:0] score_1_x470;
wire signed [DEBIT:0] score_1_x471;
wire signed [DEBIT:0] score_1_x472;
wire signed [DEBIT:0] score_1_x473;
wire signed [DEBIT:0] score_1_x474;
wire signed [DEBIT:0] score_1_x475;
wire signed [DEBIT:0] score_1_x476;
wire signed [DEBIT:0] score_1_x477;
wire signed [DEBIT:0] score_1_x478;
wire signed [DEBIT:0] score_1_x479;
wire signed [DEBIT:0] score_1_x480;
wire signed [DEBIT:0] score_1_x481;
wire signed [DEBIT:0] score_1_x482;
wire signed [DEBIT:0] score_1_x483;
wire signed [DEBIT:0] score_1_x484;
wire signed [DEBIT:0] score_1_x485;
wire signed [DEBIT:0] score_1_x486;
wire signed [DEBIT:0] score_1_x487;
wire signed [DEBIT:0] score_1_x488;
wire signed [DEBIT:0] score_1_x489;
wire signed [DEBIT:0] score_1_x490;
wire signed [DEBIT:0] score_1_x491;
wire signed [DEBIT:0] score_1_x492;
wire signed [DEBIT:0] score_1_x493;
wire signed [DEBIT:0] score_1_x494;
wire signed [DEBIT:0] score_1_x495;
wire signed [DEBIT:0] score_1_x496;
wire signed [DEBIT:0] score_1_x497;
wire signed [DEBIT:0] score_1_x498;
wire signed [DEBIT:0] score_1_x499;
wire signed [DEBIT:0] score_1_x500;
wire signed [DEBIT:0] score_1_x501;
wire signed [DEBIT:0] score_1_x502;
wire signed [DEBIT:0] score_1_x503;
wire signed [DEBIT:0] score_1_x504;
wire signed [DEBIT:0] score_1_x505;
wire signed [DEBIT:0] score_1_x506;
wire signed [DEBIT:0] score_1_x507;
wire signed [DEBIT:0] score_1_x508;
wire signed [DEBIT:0] score_1_x509;
wire signed [DEBIT:0] score_1_x510;
wire signed [DEBIT:0] score_1_x511;
wire signed [DEBIT:0] score_1_x512;
wire signed [DEBIT:0] score_1_x513;
wire signed [DEBIT:0] score_1_x514;
wire signed [DEBIT:0] score_1_x515;
wire signed [DEBIT:0] score_1_x516;
wire signed [DEBIT:0] score_1_x517;
wire signed [DEBIT:0] score_1_x518;
wire signed [DEBIT:0] score_1_x519;
wire signed [DEBIT:0] score_1_x520;
wire signed [DEBIT:0] score_1_x521;
wire signed [DEBIT:0] score_1_x522;
wire signed [DEBIT:0] score_1_x523;
wire signed [DEBIT:0] score_1_x524;
wire signed [DEBIT:0] score_1_x525;
wire signed [DEBIT:0] score_1_x526;
wire signed [DEBIT:0] score_1_x527;
wire signed [DEBIT:0] score_1_x528;
wire signed [DEBIT:0] score_1_x529;
wire signed [DEBIT:0] score_1_x530;
wire signed [DEBIT:0] score_1_x531;
wire signed [DEBIT:0] score_1_x532;
wire signed [DEBIT:0] score_1_x533;
wire signed [DEBIT:0] score_1_x534;
wire signed [DEBIT:0] score_1_x535;
wire signed [DEBIT:0] score_1_x536;
wire signed [DEBIT:0] score_1_x537;
wire signed [DEBIT:0] score_1_x538;
wire signed [DEBIT:0] score_1_x539;
wire signed [DEBIT:0] score_1_x540;
wire signed [DEBIT:0] score_1_x541;
wire signed [DEBIT:0] score_1_x542;
wire signed [DEBIT:0] score_1_x543;
wire signed [DEBIT:0] score_1_x544;
wire signed [DEBIT:0] score_1_x545;
wire signed [DEBIT:0] score_1_x546;
wire signed [DEBIT:0] score_1_x547;
wire signed [DEBIT:0] score_1_x548;
wire signed [DEBIT:0] score_1_x549;
wire signed [DEBIT:0] score_1_x550;
wire signed [DEBIT:0] score_1_x551;
wire signed [DEBIT:0] score_1_x552;
wire signed [DEBIT:0] score_1_x553;
wire signed [DEBIT:0] score_1_x554;
wire signed [DEBIT:0] score_1_x555;
wire signed [DEBIT:0] score_1_x556;
wire signed [DEBIT:0] score_1_x557;
wire signed [DEBIT:0] score_1_x558;
wire signed [DEBIT:0] score_1_x559;
wire signed [DEBIT:0] score_1_x560;
wire signed [DEBIT:0] score_1_x561;
wire signed [DEBIT:0] score_1_x562;
wire signed [DEBIT:0] score_1_x563;
wire signed [DEBIT:0] score_1_x564;
wire signed [DEBIT:0] score_1_x565;
wire signed [DEBIT:0] score_1_x566;
wire signed [DEBIT:0] score_1_x567;
wire signed [DEBIT:0] score_1_x568;
wire signed [DEBIT:0] score_1_x569;
wire signed [DEBIT:0] score_1_x570;
wire signed [DEBIT:0] score_1_x571;
wire signed [DEBIT:0] score_1_x572;
wire signed [DEBIT:0] score_1_x573;
wire signed [DEBIT:0] score_1_x574;
wire signed [DEBIT:0] score_1_x575;
wire signed [DEBIT:0] score_1_x576;
wire signed [DEBIT:0] score_1_x577;
wire signed [DEBIT:0] score_1_x578;
wire signed [DEBIT:0] score_1_x579;
wire signed [DEBIT:0] score_1_x580;
wire signed [DEBIT:0] score_1_x581;
wire signed [DEBIT:0] score_1_x582;
wire signed [DEBIT:0] score_1_x583;
wire signed [DEBIT:0] score_1_x584;
wire signed [DEBIT:0] score_1_x585;
wire signed [DEBIT:0] score_1_x586;
wire signed [DEBIT:0] score_1_x587;
wire signed [DEBIT:0] score_1_x588;
wire signed [DEBIT:0] score_1_x589;
wire signed [DEBIT:0] score_1_x590;
wire signed [DEBIT:0] score_1_x591;
wire signed [DEBIT:0] score_1_x592;
wire signed [DEBIT:0] score_1_x593;
wire signed [DEBIT:0] score_1_x594;
wire signed [DEBIT:0] score_1_x595;
wire signed [DEBIT:0] score_1_x596;
wire signed [DEBIT:0] score_1_x597;
wire signed [DEBIT:0] score_1_x598;
wire signed [DEBIT:0] score_1_x599;
wire signed [DEBIT:0] score_1_x600;
wire signed [DEBIT:0] score_1_x601;
wire signed [DEBIT:0] score_1_x602;
wire signed [DEBIT:0] score_1_x603;
wire signed [DEBIT:0] score_1_x604;
wire signed [DEBIT:0] score_1_x605;
wire signed [DEBIT:0] score_1_x606;
wire signed [DEBIT:0] score_1_x607;
wire signed [DEBIT:0] score_1_x608;
wire signed [DEBIT:0] score_1_x609;
wire signed [DEBIT:0] score_1_x610;
wire signed [DEBIT:0] score_1_x611;
wire signed [DEBIT:0] score_1_x612;
wire signed [DEBIT:0] score_1_x613;
wire signed [DEBIT:0] score_1_x614;
wire signed [DEBIT:0] score_1_x615;
wire signed [DEBIT:0] score_1_x616;
wire signed [DEBIT:0] score_1_x617;
wire signed [DEBIT:0] score_1_x618;
wire signed [DEBIT:0] score_1_x619;
wire signed [DEBIT:0] score_1_x620;
wire signed [DEBIT:0] score_1_x621;
wire signed [DEBIT:0] score_1_x622;
wire signed [DEBIT:0] score_1_x623;
wire signed [DEBIT:0] score_1_x624;
wire signed [DEBIT:0] score_1_x625;
wire signed [DEBIT:0] score_1_x626;
wire signed [DEBIT:0] score_1_x627;
wire signed [DEBIT:0] score_1_x628;
wire signed [DEBIT:0] score_1_x629;
wire signed [DEBIT:0] score_1_x630;
wire signed [DEBIT:0] score_1_x631;
wire signed [DEBIT:0] score_1_x632;
wire signed [DEBIT:0] score_1_x633;
wire signed [DEBIT:0] score_1_x634;
wire signed [DEBIT:0] score_1_x635;
wire signed [DEBIT:0] score_1_x636;
wire signed [DEBIT:0] score_1_x637;
wire signed [DEBIT:0] score_1_x638;
wire signed [DEBIT:0] score_1_x639;
wire signed [DEBIT:0] score_1_x640;
wire signed [DEBIT:0] score_1_x641;
wire signed [DEBIT:0] score_1_x642;
wire signed [DEBIT:0] score_1_x643;
wire signed [DEBIT:0] score_1_x644;
wire signed [DEBIT:0] score_1_x645;
wire signed [DEBIT:0] score_1_x646;
wire signed [DEBIT:0] score_1_x647;
wire signed [DEBIT:0] score_1_x648;
wire signed [DEBIT:0] score_1_x649;
wire signed [DEBIT:0] score_1_x650;
wire signed [DEBIT:0] score_1_x651;
wire signed [DEBIT:0] score_1_x652;
wire signed [DEBIT:0] score_1_x653;
wire signed [DEBIT:0] score_1_x654;
wire signed [DEBIT:0] score_1_x655;
wire signed [DEBIT:0] score_1_x656;
wire signed [DEBIT:0] score_1_x657;
wire signed [DEBIT:0] score_1_x658;
wire signed [DEBIT:0] score_1_x659;
wire signed [DEBIT:0] score_1_x660;
wire signed [DEBIT:0] score_1_x661;
wire signed [DEBIT:0] score_1_x662;
wire signed [DEBIT:0] score_1_x663;
wire signed [DEBIT:0] score_1_x664;
wire signed [DEBIT:0] score_1_x665;
wire signed [DEBIT:0] score_1_x666;
wire signed [DEBIT:0] score_1_x667;
wire signed [DEBIT:0] score_1_x668;
wire signed [DEBIT:0] score_1_x669;
wire signed [DEBIT:0] score_1_x670;
wire signed [DEBIT:0] score_1_x671;
wire signed [DEBIT:0] score_1_x672;
wire signed [DEBIT:0] score_1_x673;
wire signed [DEBIT:0] score_1_x674;
wire signed [DEBIT:0] score_1_x675;
wire signed [DEBIT:0] score_1_x676;
wire signed [DEBIT:0] score_1_x677;
wire signed [DEBIT:0] score_1_x678;
wire signed [DEBIT:0] score_1_x679;
wire signed [DEBIT:0] score_1_x680;
wire signed [DEBIT:0] score_1_x681;
wire signed [DEBIT:0] score_1_x682;
wire signed [DEBIT:0] score_1_x683;
wire signed [DEBIT:0] score_1_x684;
wire signed [DEBIT:0] score_1_x685;
wire signed [DEBIT:0] score_1_x686;
wire signed [DEBIT:0] score_1_x687;
wire signed [DEBIT:0] score_1_x688;
wire signed [DEBIT:0] score_1_x689;
wire signed [DEBIT:0] score_1_x690;
wire signed [DEBIT:0] score_1_x691;
wire signed [DEBIT:0] score_1_x692;
wire signed [DEBIT:0] score_1_x693;
wire signed [DEBIT:0] score_1_x694;
wire signed [DEBIT:0] score_1_x695;
wire signed [DEBIT:0] score_1_x696;
wire signed [DEBIT:0] score_1_x697;
wire signed [DEBIT:0] score_1_x698;
wire signed [DEBIT:0] score_1_x699;
wire signed [DEBIT:0] score_1_x700;
wire signed [DEBIT:0] score_1_x701;
wire signed [DEBIT:0] score_1_x702;
wire signed [DEBIT:0] score_1_x703;
wire signed [DEBIT:0] score_1_x704;
wire signed [DEBIT:0] score_1_x705;
wire signed [DEBIT:0] score_1_x706;
wire signed [DEBIT:0] score_1_x707;
wire signed [DEBIT:0] score_1_x708;
wire signed [DEBIT:0] score_1_x709;
wire signed [DEBIT:0] score_1_x710;
wire signed [DEBIT:0] score_1_x711;
wire signed [DEBIT:0] score_1_x712;
wire signed [DEBIT:0] score_1_x713;
wire signed [DEBIT:0] score_1_x714;
wire signed [DEBIT:0] score_1_x715;
wire signed [DEBIT:0] score_1_x716;
wire signed [DEBIT:0] score_1_x717;
wire signed [DEBIT:0] score_1_x718;
wire signed [DEBIT:0] score_1_x719;
wire signed [DEBIT:0] score_1_x720;
wire signed [DEBIT:0] score_1_x721;
wire signed [DEBIT:0] score_1_x722;
wire signed [DEBIT:0] score_1_x723;
wire signed [DEBIT:0] score_1_x724;
wire signed [DEBIT:0] score_1_x725;
wire signed [DEBIT:0] score_1_x726;
wire signed [DEBIT:0] score_1_x727;
wire signed [DEBIT:0] score_1_x728;
wire signed [DEBIT:0] score_1_x729;
wire signed [DEBIT:0] score_1_x730;
wire signed [DEBIT:0] score_1_x731;
wire signed [DEBIT:0] score_1_x732;
wire signed [DEBIT:0] score_1_x733;
wire signed [DEBIT:0] score_1_x734;
wire signed [DEBIT:0] score_1_x735;
wire signed [DEBIT:0] score_1_x736;
wire signed [DEBIT:0] score_1_x737;
wire signed [DEBIT:0] score_1_x738;
wire signed [DEBIT:0] score_1_x739;
wire signed [DEBIT:0] score_1_x740;
wire signed [DEBIT:0] score_1_x741;
wire signed [DEBIT:0] score_1_x742;
wire signed [DEBIT:0] score_1_x743;
wire signed [DEBIT:0] score_1_x744;
wire signed [DEBIT:0] score_1_x745;
wire signed [DEBIT:0] score_1_x746;
wire signed [DEBIT:0] score_1_x747;
wire signed [DEBIT:0] score_1_x748;
wire signed [DEBIT:0] score_1_x749;
wire signed [DEBIT:0] score_1_x750;
wire signed [DEBIT:0] score_1_x751;
wire signed [DEBIT:0] score_1_x752;
wire signed [DEBIT:0] score_1_x753;
wire signed [DEBIT:0] score_1_x754;
wire signed [DEBIT:0] score_1_x755;
wire signed [DEBIT:0] score_1_x756;
wire signed [DEBIT:0] score_1_x757;
wire signed [DEBIT:0] score_1_x758;
wire signed [DEBIT:0] score_1_x759;
wire signed [DEBIT:0] score_1_x760;
wire signed [DEBIT:0] score_1_x761;
wire signed [DEBIT:0] score_1_x762;
wire signed [DEBIT:0] score_1_x763;
wire signed [DEBIT:0] score_1_x764;
wire signed [DEBIT:0] score_1_x765;
wire signed [DEBIT:0] score_1_x766;
wire signed [DEBIT:0] score_1_x767;
wire signed [DEBIT:0] score_1_x768;
wire signed [DEBIT:0] score_1_x769;
wire signed [DEBIT:0] score_1_x770;
wire signed [DEBIT:0] score_1_x771;
wire signed [DEBIT:0] score_1_x772;
wire signed [DEBIT:0] score_1_x773;
wire signed [DEBIT:0] score_1_x774;
wire signed [DEBIT:0] score_1_x775;
wire signed [DEBIT:0] score_1_x776;
wire signed [DEBIT:0] score_1_x777;
wire signed [DEBIT:0] score_1_x778;
wire signed [DEBIT:0] score_1_x779;
wire signed [DEBIT:0] score_1_x780;
wire signed [DEBIT:0] score_1_x781;
wire signed [DEBIT:0] score_1_x782;
wire signed [DEBIT:0] score_1_x783;
wire signed [DEBIT:0] score_1_x784;
wire signed [DEBIT:0] score_2_x1;
wire signed [DEBIT:0] score_2_x2;
wire signed [DEBIT:0] score_2_x3;
wire signed [DEBIT:0] score_2_x4;
wire signed [DEBIT:0] score_2_x5;
wire signed [DEBIT:0] score_2_x6;
wire signed [DEBIT:0] score_2_x7;
wire signed [DEBIT:0] score_2_x8;
wire signed [DEBIT:0] score_2_x9;
wire signed [DEBIT:0] score_2_x10;
wire signed [DEBIT:0] score_2_x11;
wire signed [DEBIT:0] score_2_x12;
wire signed [DEBIT:0] score_2_x13;
wire signed [DEBIT:0] score_2_x14;
wire signed [DEBIT:0] score_2_x15;
wire signed [DEBIT:0] score_2_x16;
wire signed [DEBIT:0] score_2_x17;
wire signed [DEBIT:0] score_2_x18;
wire signed [DEBIT:0] score_2_x19;
wire signed [DEBIT:0] score_2_x20;
wire signed [DEBIT:0] score_2_x21;
wire signed [DEBIT:0] score_2_x22;
wire signed [DEBIT:0] score_2_x23;
wire signed [DEBIT:0] score_2_x24;
wire signed [DEBIT:0] score_2_x25;
wire signed [DEBIT:0] score_2_x26;
wire signed [DEBIT:0] score_2_x27;
wire signed [DEBIT:0] score_2_x28;
wire signed [DEBIT:0] score_2_x29;
wire signed [DEBIT:0] score_2_x30;
wire signed [DEBIT:0] score_2_x31;
wire signed [DEBIT:0] score_2_x32;
wire signed [DEBIT:0] score_2_x33;
wire signed [DEBIT:0] score_2_x34;
wire signed [DEBIT:0] score_2_x35;
wire signed [DEBIT:0] score_2_x36;
wire signed [DEBIT:0] score_2_x37;
wire signed [DEBIT:0] score_2_x38;
wire signed [DEBIT:0] score_2_x39;
wire signed [DEBIT:0] score_2_x40;
wire signed [DEBIT:0] score_2_x41;
wire signed [DEBIT:0] score_2_x42;
wire signed [DEBIT:0] score_2_x43;
wire signed [DEBIT:0] score_2_x44;
wire signed [DEBIT:0] score_2_x45;
wire signed [DEBIT:0] score_2_x46;
wire signed [DEBIT:0] score_2_x47;
wire signed [DEBIT:0] score_2_x48;
wire signed [DEBIT:0] score_2_x49;
wire signed [DEBIT:0] score_2_x50;
wire signed [DEBIT:0] score_2_x51;
wire signed [DEBIT:0] score_2_x52;
wire signed [DEBIT:0] score_2_x53;
wire signed [DEBIT:0] score_2_x54;
wire signed [DEBIT:0] score_2_x55;
wire signed [DEBIT:0] score_2_x56;
wire signed [DEBIT:0] score_2_x57;
wire signed [DEBIT:0] score_2_x58;
wire signed [DEBIT:0] score_2_x59;
wire signed [DEBIT:0] score_2_x60;
wire signed [DEBIT:0] score_2_x61;
wire signed [DEBIT:0] score_2_x62;
wire signed [DEBIT:0] score_2_x63;
wire signed [DEBIT:0] score_2_x64;
wire signed [DEBIT:0] score_2_x65;
wire signed [DEBIT:0] score_2_x66;
wire signed [DEBIT:0] score_2_x67;
wire signed [DEBIT:0] score_2_x68;
wire signed [DEBIT:0] score_2_x69;
wire signed [DEBIT:0] score_2_x70;
wire signed [DEBIT:0] score_2_x71;
wire signed [DEBIT:0] score_2_x72;
wire signed [DEBIT:0] score_2_x73;
wire signed [DEBIT:0] score_2_x74;
wire signed [DEBIT:0] score_2_x75;
wire signed [DEBIT:0] score_2_x76;
wire signed [DEBIT:0] score_2_x77;
wire signed [DEBIT:0] score_2_x78;
wire signed [DEBIT:0] score_2_x79;
wire signed [DEBIT:0] score_2_x80;
wire signed [DEBIT:0] score_2_x81;
wire signed [DEBIT:0] score_2_x82;
wire signed [DEBIT:0] score_2_x83;
wire signed [DEBIT:0] score_2_x84;
wire signed [DEBIT:0] score_2_x85;
wire signed [DEBIT:0] score_2_x86;
wire signed [DEBIT:0] score_2_x87;
wire signed [DEBIT:0] score_2_x88;
wire signed [DEBIT:0] score_2_x89;
wire signed [DEBIT:0] score_2_x90;
wire signed [DEBIT:0] score_2_x91;
wire signed [DEBIT:0] score_2_x92;
wire signed [DEBIT:0] score_2_x93;
wire signed [DEBIT:0] score_2_x94;
wire signed [DEBIT:0] score_2_x95;
wire signed [DEBIT:0] score_2_x96;
wire signed [DEBIT:0] score_2_x97;
wire signed [DEBIT:0] score_2_x98;
wire signed [DEBIT:0] score_2_x99;
wire signed [DEBIT:0] score_2_x100;
wire signed [DEBIT:0] score_2_x101;
wire signed [DEBIT:0] score_2_x102;
wire signed [DEBIT:0] score_2_x103;
wire signed [DEBIT:0] score_2_x104;
wire signed [DEBIT:0] score_2_x105;
wire signed [DEBIT:0] score_2_x106;
wire signed [DEBIT:0] score_2_x107;
wire signed [DEBIT:0] score_2_x108;
wire signed [DEBIT:0] score_2_x109;
wire signed [DEBIT:0] score_2_x110;
wire signed [DEBIT:0] score_2_x111;
wire signed [DEBIT:0] score_2_x112;
wire signed [DEBIT:0] score_2_x113;
wire signed [DEBIT:0] score_2_x114;
wire signed [DEBIT:0] score_2_x115;
wire signed [DEBIT:0] score_2_x116;
wire signed [DEBIT:0] score_2_x117;
wire signed [DEBIT:0] score_2_x118;
wire signed [DEBIT:0] score_2_x119;
wire signed [DEBIT:0] score_2_x120;
wire signed [DEBIT:0] score_2_x121;
wire signed [DEBIT:0] score_2_x122;
wire signed [DEBIT:0] score_2_x123;
wire signed [DEBIT:0] score_2_x124;
wire signed [DEBIT:0] score_2_x125;
wire signed [DEBIT:0] score_2_x126;
wire signed [DEBIT:0] score_2_x127;
wire signed [DEBIT:0] score_2_x128;
wire signed [DEBIT:0] score_2_x129;
wire signed [DEBIT:0] score_2_x130;
wire signed [DEBIT:0] score_2_x131;
wire signed [DEBIT:0] score_2_x132;
wire signed [DEBIT:0] score_2_x133;
wire signed [DEBIT:0] score_2_x134;
wire signed [DEBIT:0] score_2_x135;
wire signed [DEBIT:0] score_2_x136;
wire signed [DEBIT:0] score_2_x137;
wire signed [DEBIT:0] score_2_x138;
wire signed [DEBIT:0] score_2_x139;
wire signed [DEBIT:0] score_2_x140;
wire signed [DEBIT:0] score_2_x141;
wire signed [DEBIT:0] score_2_x142;
wire signed [DEBIT:0] score_2_x143;
wire signed [DEBIT:0] score_2_x144;
wire signed [DEBIT:0] score_2_x145;
wire signed [DEBIT:0] score_2_x146;
wire signed [DEBIT:0] score_2_x147;
wire signed [DEBIT:0] score_2_x148;
wire signed [DEBIT:0] score_2_x149;
wire signed [DEBIT:0] score_2_x150;
wire signed [DEBIT:0] score_2_x151;
wire signed [DEBIT:0] score_2_x152;
wire signed [DEBIT:0] score_2_x153;
wire signed [DEBIT:0] score_2_x154;
wire signed [DEBIT:0] score_2_x155;
wire signed [DEBIT:0] score_2_x156;
wire signed [DEBIT:0] score_2_x157;
wire signed [DEBIT:0] score_2_x158;
wire signed [DEBIT:0] score_2_x159;
wire signed [DEBIT:0] score_2_x160;
wire signed [DEBIT:0] score_2_x161;
wire signed [DEBIT:0] score_2_x162;
wire signed [DEBIT:0] score_2_x163;
wire signed [DEBIT:0] score_2_x164;
wire signed [DEBIT:0] score_2_x165;
wire signed [DEBIT:0] score_2_x166;
wire signed [DEBIT:0] score_2_x167;
wire signed [DEBIT:0] score_2_x168;
wire signed [DEBIT:0] score_2_x169;
wire signed [DEBIT:0] score_2_x170;
wire signed [DEBIT:0] score_2_x171;
wire signed [DEBIT:0] score_2_x172;
wire signed [DEBIT:0] score_2_x173;
wire signed [DEBIT:0] score_2_x174;
wire signed [DEBIT:0] score_2_x175;
wire signed [DEBIT:0] score_2_x176;
wire signed [DEBIT:0] score_2_x177;
wire signed [DEBIT:0] score_2_x178;
wire signed [DEBIT:0] score_2_x179;
wire signed [DEBIT:0] score_2_x180;
wire signed [DEBIT:0] score_2_x181;
wire signed [DEBIT:0] score_2_x182;
wire signed [DEBIT:0] score_2_x183;
wire signed [DEBIT:0] score_2_x184;
wire signed [DEBIT:0] score_2_x185;
wire signed [DEBIT:0] score_2_x186;
wire signed [DEBIT:0] score_2_x187;
wire signed [DEBIT:0] score_2_x188;
wire signed [DEBIT:0] score_2_x189;
wire signed [DEBIT:0] score_2_x190;
wire signed [DEBIT:0] score_2_x191;
wire signed [DEBIT:0] score_2_x192;
wire signed [DEBIT:0] score_2_x193;
wire signed [DEBIT:0] score_2_x194;
wire signed [DEBIT:0] score_2_x195;
wire signed [DEBIT:0] score_2_x196;
wire signed [DEBIT:0] score_2_x197;
wire signed [DEBIT:0] score_2_x198;
wire signed [DEBIT:0] score_2_x199;
wire signed [DEBIT:0] score_2_x200;
wire signed [DEBIT:0] score_2_x201;
wire signed [DEBIT:0] score_2_x202;
wire signed [DEBIT:0] score_2_x203;
wire signed [DEBIT:0] score_2_x204;
wire signed [DEBIT:0] score_2_x205;
wire signed [DEBIT:0] score_2_x206;
wire signed [DEBIT:0] score_2_x207;
wire signed [DEBIT:0] score_2_x208;
wire signed [DEBIT:0] score_2_x209;
wire signed [DEBIT:0] score_2_x210;
wire signed [DEBIT:0] score_2_x211;
wire signed [DEBIT:0] score_2_x212;
wire signed [DEBIT:0] score_2_x213;
wire signed [DEBIT:0] score_2_x214;
wire signed [DEBIT:0] score_2_x215;
wire signed [DEBIT:0] score_2_x216;
wire signed [DEBIT:0] score_2_x217;
wire signed [DEBIT:0] score_2_x218;
wire signed [DEBIT:0] score_2_x219;
wire signed [DEBIT:0] score_2_x220;
wire signed [DEBIT:0] score_2_x221;
wire signed [DEBIT:0] score_2_x222;
wire signed [DEBIT:0] score_2_x223;
wire signed [DEBIT:0] score_2_x224;
wire signed [DEBIT:0] score_2_x225;
wire signed [DEBIT:0] score_2_x226;
wire signed [DEBIT:0] score_2_x227;
wire signed [DEBIT:0] score_2_x228;
wire signed [DEBIT:0] score_2_x229;
wire signed [DEBIT:0] score_2_x230;
wire signed [DEBIT:0] score_2_x231;
wire signed [DEBIT:0] score_2_x232;
wire signed [DEBIT:0] score_2_x233;
wire signed [DEBIT:0] score_2_x234;
wire signed [DEBIT:0] score_2_x235;
wire signed [DEBIT:0] score_2_x236;
wire signed [DEBIT:0] score_2_x237;
wire signed [DEBIT:0] score_2_x238;
wire signed [DEBIT:0] score_2_x239;
wire signed [DEBIT:0] score_2_x240;
wire signed [DEBIT:0] score_2_x241;
wire signed [DEBIT:0] score_2_x242;
wire signed [DEBIT:0] score_2_x243;
wire signed [DEBIT:0] score_2_x244;
wire signed [DEBIT:0] score_2_x245;
wire signed [DEBIT:0] score_2_x246;
wire signed [DEBIT:0] score_2_x247;
wire signed [DEBIT:0] score_2_x248;
wire signed [DEBIT:0] score_2_x249;
wire signed [DEBIT:0] score_2_x250;
wire signed [DEBIT:0] score_2_x251;
wire signed [DEBIT:0] score_2_x252;
wire signed [DEBIT:0] score_2_x253;
wire signed [DEBIT:0] score_2_x254;
wire signed [DEBIT:0] score_2_x255;
wire signed [DEBIT:0] score_2_x256;
wire signed [DEBIT:0] score_2_x257;
wire signed [DEBIT:0] score_2_x258;
wire signed [DEBIT:0] score_2_x259;
wire signed [DEBIT:0] score_2_x260;
wire signed [DEBIT:0] score_2_x261;
wire signed [DEBIT:0] score_2_x262;
wire signed [DEBIT:0] score_2_x263;
wire signed [DEBIT:0] score_2_x264;
wire signed [DEBIT:0] score_2_x265;
wire signed [DEBIT:0] score_2_x266;
wire signed [DEBIT:0] score_2_x267;
wire signed [DEBIT:0] score_2_x268;
wire signed [DEBIT:0] score_2_x269;
wire signed [DEBIT:0] score_2_x270;
wire signed [DEBIT:0] score_2_x271;
wire signed [DEBIT:0] score_2_x272;
wire signed [DEBIT:0] score_2_x273;
wire signed [DEBIT:0] score_2_x274;
wire signed [DEBIT:0] score_2_x275;
wire signed [DEBIT:0] score_2_x276;
wire signed [DEBIT:0] score_2_x277;
wire signed [DEBIT:0] score_2_x278;
wire signed [DEBIT:0] score_2_x279;
wire signed [DEBIT:0] score_2_x280;
wire signed [DEBIT:0] score_2_x281;
wire signed [DEBIT:0] score_2_x282;
wire signed [DEBIT:0] score_2_x283;
wire signed [DEBIT:0] score_2_x284;
wire signed [DEBIT:0] score_2_x285;
wire signed [DEBIT:0] score_2_x286;
wire signed [DEBIT:0] score_2_x287;
wire signed [DEBIT:0] score_2_x288;
wire signed [DEBIT:0] score_2_x289;
wire signed [DEBIT:0] score_2_x290;
wire signed [DEBIT:0] score_2_x291;
wire signed [DEBIT:0] score_2_x292;
wire signed [DEBIT:0] score_2_x293;
wire signed [DEBIT:0] score_2_x294;
wire signed [DEBIT:0] score_2_x295;
wire signed [DEBIT:0] score_2_x296;
wire signed [DEBIT:0] score_2_x297;
wire signed [DEBIT:0] score_2_x298;
wire signed [DEBIT:0] score_2_x299;
wire signed [DEBIT:0] score_2_x300;
wire signed [DEBIT:0] score_2_x301;
wire signed [DEBIT:0] score_2_x302;
wire signed [DEBIT:0] score_2_x303;
wire signed [DEBIT:0] score_2_x304;
wire signed [DEBIT:0] score_2_x305;
wire signed [DEBIT:0] score_2_x306;
wire signed [DEBIT:0] score_2_x307;
wire signed [DEBIT:0] score_2_x308;
wire signed [DEBIT:0] score_2_x309;
wire signed [DEBIT:0] score_2_x310;
wire signed [DEBIT:0] score_2_x311;
wire signed [DEBIT:0] score_2_x312;
wire signed [DEBIT:0] score_2_x313;
wire signed [DEBIT:0] score_2_x314;
wire signed [DEBIT:0] score_2_x315;
wire signed [DEBIT:0] score_2_x316;
wire signed [DEBIT:0] score_2_x317;
wire signed [DEBIT:0] score_2_x318;
wire signed [DEBIT:0] score_2_x319;
wire signed [DEBIT:0] score_2_x320;
wire signed [DEBIT:0] score_2_x321;
wire signed [DEBIT:0] score_2_x322;
wire signed [DEBIT:0] score_2_x323;
wire signed [DEBIT:0] score_2_x324;
wire signed [DEBIT:0] score_2_x325;
wire signed [DEBIT:0] score_2_x326;
wire signed [DEBIT:0] score_2_x327;
wire signed [DEBIT:0] score_2_x328;
wire signed [DEBIT:0] score_2_x329;
wire signed [DEBIT:0] score_2_x330;
wire signed [DEBIT:0] score_2_x331;
wire signed [DEBIT:0] score_2_x332;
wire signed [DEBIT:0] score_2_x333;
wire signed [DEBIT:0] score_2_x334;
wire signed [DEBIT:0] score_2_x335;
wire signed [DEBIT:0] score_2_x336;
wire signed [DEBIT:0] score_2_x337;
wire signed [DEBIT:0] score_2_x338;
wire signed [DEBIT:0] score_2_x339;
wire signed [DEBIT:0] score_2_x340;
wire signed [DEBIT:0] score_2_x341;
wire signed [DEBIT:0] score_2_x342;
wire signed [DEBIT:0] score_2_x343;
wire signed [DEBIT:0] score_2_x344;
wire signed [DEBIT:0] score_2_x345;
wire signed [DEBIT:0] score_2_x346;
wire signed [DEBIT:0] score_2_x347;
wire signed [DEBIT:0] score_2_x348;
wire signed [DEBIT:0] score_2_x349;
wire signed [DEBIT:0] score_2_x350;
wire signed [DEBIT:0] score_2_x351;
wire signed [DEBIT:0] score_2_x352;
wire signed [DEBIT:0] score_2_x353;
wire signed [DEBIT:0] score_2_x354;
wire signed [DEBIT:0] score_2_x355;
wire signed [DEBIT:0] score_2_x356;
wire signed [DEBIT:0] score_2_x357;
wire signed [DEBIT:0] score_2_x358;
wire signed [DEBIT:0] score_2_x359;
wire signed [DEBIT:0] score_2_x360;
wire signed [DEBIT:0] score_2_x361;
wire signed [DEBIT:0] score_2_x362;
wire signed [DEBIT:0] score_2_x363;
wire signed [DEBIT:0] score_2_x364;
wire signed [DEBIT:0] score_2_x365;
wire signed [DEBIT:0] score_2_x366;
wire signed [DEBIT:0] score_2_x367;
wire signed [DEBIT:0] score_2_x368;
wire signed [DEBIT:0] score_2_x369;
wire signed [DEBIT:0] score_2_x370;
wire signed [DEBIT:0] score_2_x371;
wire signed [DEBIT:0] score_2_x372;
wire signed [DEBIT:0] score_2_x373;
wire signed [DEBIT:0] score_2_x374;
wire signed [DEBIT:0] score_2_x375;
wire signed [DEBIT:0] score_2_x376;
wire signed [DEBIT:0] score_2_x377;
wire signed [DEBIT:0] score_2_x378;
wire signed [DEBIT:0] score_2_x379;
wire signed [DEBIT:0] score_2_x380;
wire signed [DEBIT:0] score_2_x381;
wire signed [DEBIT:0] score_2_x382;
wire signed [DEBIT:0] score_2_x383;
wire signed [DEBIT:0] score_2_x384;
wire signed [DEBIT:0] score_2_x385;
wire signed [DEBIT:0] score_2_x386;
wire signed [DEBIT:0] score_2_x387;
wire signed [DEBIT:0] score_2_x388;
wire signed [DEBIT:0] score_2_x389;
wire signed [DEBIT:0] score_2_x390;
wire signed [DEBIT:0] score_2_x391;
wire signed [DEBIT:0] score_2_x392;
wire signed [DEBIT:0] score_2_x393;
wire signed [DEBIT:0] score_2_x394;
wire signed [DEBIT:0] score_2_x395;
wire signed [DEBIT:0] score_2_x396;
wire signed [DEBIT:0] score_2_x397;
wire signed [DEBIT:0] score_2_x398;
wire signed [DEBIT:0] score_2_x399;
wire signed [DEBIT:0] score_2_x400;
wire signed [DEBIT:0] score_2_x401;
wire signed [DEBIT:0] score_2_x402;
wire signed [DEBIT:0] score_2_x403;
wire signed [DEBIT:0] score_2_x404;
wire signed [DEBIT:0] score_2_x405;
wire signed [DEBIT:0] score_2_x406;
wire signed [DEBIT:0] score_2_x407;
wire signed [DEBIT:0] score_2_x408;
wire signed [DEBIT:0] score_2_x409;
wire signed [DEBIT:0] score_2_x410;
wire signed [DEBIT:0] score_2_x411;
wire signed [DEBIT:0] score_2_x412;
wire signed [DEBIT:0] score_2_x413;
wire signed [DEBIT:0] score_2_x414;
wire signed [DEBIT:0] score_2_x415;
wire signed [DEBIT:0] score_2_x416;
wire signed [DEBIT:0] score_2_x417;
wire signed [DEBIT:0] score_2_x418;
wire signed [DEBIT:0] score_2_x419;
wire signed [DEBIT:0] score_2_x420;
wire signed [DEBIT:0] score_2_x421;
wire signed [DEBIT:0] score_2_x422;
wire signed [DEBIT:0] score_2_x423;
wire signed [DEBIT:0] score_2_x424;
wire signed [DEBIT:0] score_2_x425;
wire signed [DEBIT:0] score_2_x426;
wire signed [DEBIT:0] score_2_x427;
wire signed [DEBIT:0] score_2_x428;
wire signed [DEBIT:0] score_2_x429;
wire signed [DEBIT:0] score_2_x430;
wire signed [DEBIT:0] score_2_x431;
wire signed [DEBIT:0] score_2_x432;
wire signed [DEBIT:0] score_2_x433;
wire signed [DEBIT:0] score_2_x434;
wire signed [DEBIT:0] score_2_x435;
wire signed [DEBIT:0] score_2_x436;
wire signed [DEBIT:0] score_2_x437;
wire signed [DEBIT:0] score_2_x438;
wire signed [DEBIT:0] score_2_x439;
wire signed [DEBIT:0] score_2_x440;
wire signed [DEBIT:0] score_2_x441;
wire signed [DEBIT:0] score_2_x442;
wire signed [DEBIT:0] score_2_x443;
wire signed [DEBIT:0] score_2_x444;
wire signed [DEBIT:0] score_2_x445;
wire signed [DEBIT:0] score_2_x446;
wire signed [DEBIT:0] score_2_x447;
wire signed [DEBIT:0] score_2_x448;
wire signed [DEBIT:0] score_2_x449;
wire signed [DEBIT:0] score_2_x450;
wire signed [DEBIT:0] score_2_x451;
wire signed [DEBIT:0] score_2_x452;
wire signed [DEBIT:0] score_2_x453;
wire signed [DEBIT:0] score_2_x454;
wire signed [DEBIT:0] score_2_x455;
wire signed [DEBIT:0] score_2_x456;
wire signed [DEBIT:0] score_2_x457;
wire signed [DEBIT:0] score_2_x458;
wire signed [DEBIT:0] score_2_x459;
wire signed [DEBIT:0] score_2_x460;
wire signed [DEBIT:0] score_2_x461;
wire signed [DEBIT:0] score_2_x462;
wire signed [DEBIT:0] score_2_x463;
wire signed [DEBIT:0] score_2_x464;
wire signed [DEBIT:0] score_2_x465;
wire signed [DEBIT:0] score_2_x466;
wire signed [DEBIT:0] score_2_x467;
wire signed [DEBIT:0] score_2_x468;
wire signed [DEBIT:0] score_2_x469;
wire signed [DEBIT:0] score_2_x470;
wire signed [DEBIT:0] score_2_x471;
wire signed [DEBIT:0] score_2_x472;
wire signed [DEBIT:0] score_2_x473;
wire signed [DEBIT:0] score_2_x474;
wire signed [DEBIT:0] score_2_x475;
wire signed [DEBIT:0] score_2_x476;
wire signed [DEBIT:0] score_2_x477;
wire signed [DEBIT:0] score_2_x478;
wire signed [DEBIT:0] score_2_x479;
wire signed [DEBIT:0] score_2_x480;
wire signed [DEBIT:0] score_2_x481;
wire signed [DEBIT:0] score_2_x482;
wire signed [DEBIT:0] score_2_x483;
wire signed [DEBIT:0] score_2_x484;
wire signed [DEBIT:0] score_2_x485;
wire signed [DEBIT:0] score_2_x486;
wire signed [DEBIT:0] score_2_x487;
wire signed [DEBIT:0] score_2_x488;
wire signed [DEBIT:0] score_2_x489;
wire signed [DEBIT:0] score_2_x490;
wire signed [DEBIT:0] score_2_x491;
wire signed [DEBIT:0] score_2_x492;
wire signed [DEBIT:0] score_2_x493;
wire signed [DEBIT:0] score_2_x494;
wire signed [DEBIT:0] score_2_x495;
wire signed [DEBIT:0] score_2_x496;
wire signed [DEBIT:0] score_2_x497;
wire signed [DEBIT:0] score_2_x498;
wire signed [DEBIT:0] score_2_x499;
wire signed [DEBIT:0] score_2_x500;
wire signed [DEBIT:0] score_2_x501;
wire signed [DEBIT:0] score_2_x502;
wire signed [DEBIT:0] score_2_x503;
wire signed [DEBIT:0] score_2_x504;
wire signed [DEBIT:0] score_2_x505;
wire signed [DEBIT:0] score_2_x506;
wire signed [DEBIT:0] score_2_x507;
wire signed [DEBIT:0] score_2_x508;
wire signed [DEBIT:0] score_2_x509;
wire signed [DEBIT:0] score_2_x510;
wire signed [DEBIT:0] score_2_x511;
wire signed [DEBIT:0] score_2_x512;
wire signed [DEBIT:0] score_2_x513;
wire signed [DEBIT:0] score_2_x514;
wire signed [DEBIT:0] score_2_x515;
wire signed [DEBIT:0] score_2_x516;
wire signed [DEBIT:0] score_2_x517;
wire signed [DEBIT:0] score_2_x518;
wire signed [DEBIT:0] score_2_x519;
wire signed [DEBIT:0] score_2_x520;
wire signed [DEBIT:0] score_2_x521;
wire signed [DEBIT:0] score_2_x522;
wire signed [DEBIT:0] score_2_x523;
wire signed [DEBIT:0] score_2_x524;
wire signed [DEBIT:0] score_2_x525;
wire signed [DEBIT:0] score_2_x526;
wire signed [DEBIT:0] score_2_x527;
wire signed [DEBIT:0] score_2_x528;
wire signed [DEBIT:0] score_2_x529;
wire signed [DEBIT:0] score_2_x530;
wire signed [DEBIT:0] score_2_x531;
wire signed [DEBIT:0] score_2_x532;
wire signed [DEBIT:0] score_2_x533;
wire signed [DEBIT:0] score_2_x534;
wire signed [DEBIT:0] score_2_x535;
wire signed [DEBIT:0] score_2_x536;
wire signed [DEBIT:0] score_2_x537;
wire signed [DEBIT:0] score_2_x538;
wire signed [DEBIT:0] score_2_x539;
wire signed [DEBIT:0] score_2_x540;
wire signed [DEBIT:0] score_2_x541;
wire signed [DEBIT:0] score_2_x542;
wire signed [DEBIT:0] score_2_x543;
wire signed [DEBIT:0] score_2_x544;
wire signed [DEBIT:0] score_2_x545;
wire signed [DEBIT:0] score_2_x546;
wire signed [DEBIT:0] score_2_x547;
wire signed [DEBIT:0] score_2_x548;
wire signed [DEBIT:0] score_2_x549;
wire signed [DEBIT:0] score_2_x550;
wire signed [DEBIT:0] score_2_x551;
wire signed [DEBIT:0] score_2_x552;
wire signed [DEBIT:0] score_2_x553;
wire signed [DEBIT:0] score_2_x554;
wire signed [DEBIT:0] score_2_x555;
wire signed [DEBIT:0] score_2_x556;
wire signed [DEBIT:0] score_2_x557;
wire signed [DEBIT:0] score_2_x558;
wire signed [DEBIT:0] score_2_x559;
wire signed [DEBIT:0] score_2_x560;
wire signed [DEBIT:0] score_2_x561;
wire signed [DEBIT:0] score_2_x562;
wire signed [DEBIT:0] score_2_x563;
wire signed [DEBIT:0] score_2_x564;
wire signed [DEBIT:0] score_2_x565;
wire signed [DEBIT:0] score_2_x566;
wire signed [DEBIT:0] score_2_x567;
wire signed [DEBIT:0] score_2_x568;
wire signed [DEBIT:0] score_2_x569;
wire signed [DEBIT:0] score_2_x570;
wire signed [DEBIT:0] score_2_x571;
wire signed [DEBIT:0] score_2_x572;
wire signed [DEBIT:0] score_2_x573;
wire signed [DEBIT:0] score_2_x574;
wire signed [DEBIT:0] score_2_x575;
wire signed [DEBIT:0] score_2_x576;
wire signed [DEBIT:0] score_2_x577;
wire signed [DEBIT:0] score_2_x578;
wire signed [DEBIT:0] score_2_x579;
wire signed [DEBIT:0] score_2_x580;
wire signed [DEBIT:0] score_2_x581;
wire signed [DEBIT:0] score_2_x582;
wire signed [DEBIT:0] score_2_x583;
wire signed [DEBIT:0] score_2_x584;
wire signed [DEBIT:0] score_2_x585;
wire signed [DEBIT:0] score_2_x586;
wire signed [DEBIT:0] score_2_x587;
wire signed [DEBIT:0] score_2_x588;
wire signed [DEBIT:0] score_2_x589;
wire signed [DEBIT:0] score_2_x590;
wire signed [DEBIT:0] score_2_x591;
wire signed [DEBIT:0] score_2_x592;
wire signed [DEBIT:0] score_2_x593;
wire signed [DEBIT:0] score_2_x594;
wire signed [DEBIT:0] score_2_x595;
wire signed [DEBIT:0] score_2_x596;
wire signed [DEBIT:0] score_2_x597;
wire signed [DEBIT:0] score_2_x598;
wire signed [DEBIT:0] score_2_x599;
wire signed [DEBIT:0] score_2_x600;
wire signed [DEBIT:0] score_2_x601;
wire signed [DEBIT:0] score_2_x602;
wire signed [DEBIT:0] score_2_x603;
wire signed [DEBIT:0] score_2_x604;
wire signed [DEBIT:0] score_2_x605;
wire signed [DEBIT:0] score_2_x606;
wire signed [DEBIT:0] score_2_x607;
wire signed [DEBIT:0] score_2_x608;
wire signed [DEBIT:0] score_2_x609;
wire signed [DEBIT:0] score_2_x610;
wire signed [DEBIT:0] score_2_x611;
wire signed [DEBIT:0] score_2_x612;
wire signed [DEBIT:0] score_2_x613;
wire signed [DEBIT:0] score_2_x614;
wire signed [DEBIT:0] score_2_x615;
wire signed [DEBIT:0] score_2_x616;
wire signed [DEBIT:0] score_2_x617;
wire signed [DEBIT:0] score_2_x618;
wire signed [DEBIT:0] score_2_x619;
wire signed [DEBIT:0] score_2_x620;
wire signed [DEBIT:0] score_2_x621;
wire signed [DEBIT:0] score_2_x622;
wire signed [DEBIT:0] score_2_x623;
wire signed [DEBIT:0] score_2_x624;
wire signed [DEBIT:0] score_2_x625;
wire signed [DEBIT:0] score_2_x626;
wire signed [DEBIT:0] score_2_x627;
wire signed [DEBIT:0] score_2_x628;
wire signed [DEBIT:0] score_2_x629;
wire signed [DEBIT:0] score_2_x630;
wire signed [DEBIT:0] score_2_x631;
wire signed [DEBIT:0] score_2_x632;
wire signed [DEBIT:0] score_2_x633;
wire signed [DEBIT:0] score_2_x634;
wire signed [DEBIT:0] score_2_x635;
wire signed [DEBIT:0] score_2_x636;
wire signed [DEBIT:0] score_2_x637;
wire signed [DEBIT:0] score_2_x638;
wire signed [DEBIT:0] score_2_x639;
wire signed [DEBIT:0] score_2_x640;
wire signed [DEBIT:0] score_2_x641;
wire signed [DEBIT:0] score_2_x642;
wire signed [DEBIT:0] score_2_x643;
wire signed [DEBIT:0] score_2_x644;
wire signed [DEBIT:0] score_2_x645;
wire signed [DEBIT:0] score_2_x646;
wire signed [DEBIT:0] score_2_x647;
wire signed [DEBIT:0] score_2_x648;
wire signed [DEBIT:0] score_2_x649;
wire signed [DEBIT:0] score_2_x650;
wire signed [DEBIT:0] score_2_x651;
wire signed [DEBIT:0] score_2_x652;
wire signed [DEBIT:0] score_2_x653;
wire signed [DEBIT:0] score_2_x654;
wire signed [DEBIT:0] score_2_x655;
wire signed [DEBIT:0] score_2_x656;
wire signed [DEBIT:0] score_2_x657;
wire signed [DEBIT:0] score_2_x658;
wire signed [DEBIT:0] score_2_x659;
wire signed [DEBIT:0] score_2_x660;
wire signed [DEBIT:0] score_2_x661;
wire signed [DEBIT:0] score_2_x662;
wire signed [DEBIT:0] score_2_x663;
wire signed [DEBIT:0] score_2_x664;
wire signed [DEBIT:0] score_2_x665;
wire signed [DEBIT:0] score_2_x666;
wire signed [DEBIT:0] score_2_x667;
wire signed [DEBIT:0] score_2_x668;
wire signed [DEBIT:0] score_2_x669;
wire signed [DEBIT:0] score_2_x670;
wire signed [DEBIT:0] score_2_x671;
wire signed [DEBIT:0] score_2_x672;
wire signed [DEBIT:0] score_2_x673;
wire signed [DEBIT:0] score_2_x674;
wire signed [DEBIT:0] score_2_x675;
wire signed [DEBIT:0] score_2_x676;
wire signed [DEBIT:0] score_2_x677;
wire signed [DEBIT:0] score_2_x678;
wire signed [DEBIT:0] score_2_x679;
wire signed [DEBIT:0] score_2_x680;
wire signed [DEBIT:0] score_2_x681;
wire signed [DEBIT:0] score_2_x682;
wire signed [DEBIT:0] score_2_x683;
wire signed [DEBIT:0] score_2_x684;
wire signed [DEBIT:0] score_2_x685;
wire signed [DEBIT:0] score_2_x686;
wire signed [DEBIT:0] score_2_x687;
wire signed [DEBIT:0] score_2_x688;
wire signed [DEBIT:0] score_2_x689;
wire signed [DEBIT:0] score_2_x690;
wire signed [DEBIT:0] score_2_x691;
wire signed [DEBIT:0] score_2_x692;
wire signed [DEBIT:0] score_2_x693;
wire signed [DEBIT:0] score_2_x694;
wire signed [DEBIT:0] score_2_x695;
wire signed [DEBIT:0] score_2_x696;
wire signed [DEBIT:0] score_2_x697;
wire signed [DEBIT:0] score_2_x698;
wire signed [DEBIT:0] score_2_x699;
wire signed [DEBIT:0] score_2_x700;
wire signed [DEBIT:0] score_2_x701;
wire signed [DEBIT:0] score_2_x702;
wire signed [DEBIT:0] score_2_x703;
wire signed [DEBIT:0] score_2_x704;
wire signed [DEBIT:0] score_2_x705;
wire signed [DEBIT:0] score_2_x706;
wire signed [DEBIT:0] score_2_x707;
wire signed [DEBIT:0] score_2_x708;
wire signed [DEBIT:0] score_2_x709;
wire signed [DEBIT:0] score_2_x710;
wire signed [DEBIT:0] score_2_x711;
wire signed [DEBIT:0] score_2_x712;
wire signed [DEBIT:0] score_2_x713;
wire signed [DEBIT:0] score_2_x714;
wire signed [DEBIT:0] score_2_x715;
wire signed [DEBIT:0] score_2_x716;
wire signed [DEBIT:0] score_2_x717;
wire signed [DEBIT:0] score_2_x718;
wire signed [DEBIT:0] score_2_x719;
wire signed [DEBIT:0] score_2_x720;
wire signed [DEBIT:0] score_2_x721;
wire signed [DEBIT:0] score_2_x722;
wire signed [DEBIT:0] score_2_x723;
wire signed [DEBIT:0] score_2_x724;
wire signed [DEBIT:0] score_2_x725;
wire signed [DEBIT:0] score_2_x726;
wire signed [DEBIT:0] score_2_x727;
wire signed [DEBIT:0] score_2_x728;
wire signed [DEBIT:0] score_2_x729;
wire signed [DEBIT:0] score_2_x730;
wire signed [DEBIT:0] score_2_x731;
wire signed [DEBIT:0] score_2_x732;
wire signed [DEBIT:0] score_2_x733;
wire signed [DEBIT:0] score_2_x734;
wire signed [DEBIT:0] score_2_x735;
wire signed [DEBIT:0] score_2_x736;
wire signed [DEBIT:0] score_2_x737;
wire signed [DEBIT:0] score_2_x738;
wire signed [DEBIT:0] score_2_x739;
wire signed [DEBIT:0] score_2_x740;
wire signed [DEBIT:0] score_2_x741;
wire signed [DEBIT:0] score_2_x742;
wire signed [DEBIT:0] score_2_x743;
wire signed [DEBIT:0] score_2_x744;
wire signed [DEBIT:0] score_2_x745;
wire signed [DEBIT:0] score_2_x746;
wire signed [DEBIT:0] score_2_x747;
wire signed [DEBIT:0] score_2_x748;
wire signed [DEBIT:0] score_2_x749;
wire signed [DEBIT:0] score_2_x750;
wire signed [DEBIT:0] score_2_x751;
wire signed [DEBIT:0] score_2_x752;
wire signed [DEBIT:0] score_2_x753;
wire signed [DEBIT:0] score_2_x754;
wire signed [DEBIT:0] score_2_x755;
wire signed [DEBIT:0] score_2_x756;
wire signed [DEBIT:0] score_2_x757;
wire signed [DEBIT:0] score_2_x758;
wire signed [DEBIT:0] score_2_x759;
wire signed [DEBIT:0] score_2_x760;
wire signed [DEBIT:0] score_2_x761;
wire signed [DEBIT:0] score_2_x762;
wire signed [DEBIT:0] score_2_x763;
wire signed [DEBIT:0] score_2_x764;
wire signed [DEBIT:0] score_2_x765;
wire signed [DEBIT:0] score_2_x766;
wire signed [DEBIT:0] score_2_x767;
wire signed [DEBIT:0] score_2_x768;
wire signed [DEBIT:0] score_2_x769;
wire signed [DEBIT:0] score_2_x770;
wire signed [DEBIT:0] score_2_x771;
wire signed [DEBIT:0] score_2_x772;
wire signed [DEBIT:0] score_2_x773;
wire signed [DEBIT:0] score_2_x774;
wire signed [DEBIT:0] score_2_x775;
wire signed [DEBIT:0] score_2_x776;
wire signed [DEBIT:0] score_2_x777;
wire signed [DEBIT:0] score_2_x778;
wire signed [DEBIT:0] score_2_x779;
wire signed [DEBIT:0] score_2_x780;
wire signed [DEBIT:0] score_2_x781;
wire signed [DEBIT:0] score_2_x782;
wire signed [DEBIT:0] score_2_x783;
wire signed [DEBIT:0] score_2_x784;
wire signed [DEBIT:0] score_3_x1;
wire signed [DEBIT:0] score_3_x2;
wire signed [DEBIT:0] score_3_x3;
wire signed [DEBIT:0] score_3_x4;
wire signed [DEBIT:0] score_3_x5;
wire signed [DEBIT:0] score_3_x6;
wire signed [DEBIT:0] score_3_x7;
wire signed [DEBIT:0] score_3_x8;
wire signed [DEBIT:0] score_3_x9;
wire signed [DEBIT:0] score_3_x10;
wire signed [DEBIT:0] score_3_x11;
wire signed [DEBIT:0] score_3_x12;
wire signed [DEBIT:0] score_3_x13;
wire signed [DEBIT:0] score_3_x14;
wire signed [DEBIT:0] score_3_x15;
wire signed [DEBIT:0] score_3_x16;
wire signed [DEBIT:0] score_3_x17;
wire signed [DEBIT:0] score_3_x18;
wire signed [DEBIT:0] score_3_x19;
wire signed [DEBIT:0] score_3_x20;
wire signed [DEBIT:0] score_3_x21;
wire signed [DEBIT:0] score_3_x22;
wire signed [DEBIT:0] score_3_x23;
wire signed [DEBIT:0] score_3_x24;
wire signed [DEBIT:0] score_3_x25;
wire signed [DEBIT:0] score_3_x26;
wire signed [DEBIT:0] score_3_x27;
wire signed [DEBIT:0] score_3_x28;
wire signed [DEBIT:0] score_3_x29;
wire signed [DEBIT:0] score_3_x30;
wire signed [DEBIT:0] score_3_x31;
wire signed [DEBIT:0] score_3_x32;
wire signed [DEBIT:0] score_3_x33;
wire signed [DEBIT:0] score_3_x34;
wire signed [DEBIT:0] score_3_x35;
wire signed [DEBIT:0] score_3_x36;
wire signed [DEBIT:0] score_3_x37;
wire signed [DEBIT:0] score_3_x38;
wire signed [DEBIT:0] score_3_x39;
wire signed [DEBIT:0] score_3_x40;
wire signed [DEBIT:0] score_3_x41;
wire signed [DEBIT:0] score_3_x42;
wire signed [DEBIT:0] score_3_x43;
wire signed [DEBIT:0] score_3_x44;
wire signed [DEBIT:0] score_3_x45;
wire signed [DEBIT:0] score_3_x46;
wire signed [DEBIT:0] score_3_x47;
wire signed [DEBIT:0] score_3_x48;
wire signed [DEBIT:0] score_3_x49;
wire signed [DEBIT:0] score_3_x50;
wire signed [DEBIT:0] score_3_x51;
wire signed [DEBIT:0] score_3_x52;
wire signed [DEBIT:0] score_3_x53;
wire signed [DEBIT:0] score_3_x54;
wire signed [DEBIT:0] score_3_x55;
wire signed [DEBIT:0] score_3_x56;
wire signed [DEBIT:0] score_3_x57;
wire signed [DEBIT:0] score_3_x58;
wire signed [DEBIT:0] score_3_x59;
wire signed [DEBIT:0] score_3_x60;
wire signed [DEBIT:0] score_3_x61;
wire signed [DEBIT:0] score_3_x62;
wire signed [DEBIT:0] score_3_x63;
wire signed [DEBIT:0] score_3_x64;
wire signed [DEBIT:0] score_3_x65;
wire signed [DEBIT:0] score_3_x66;
wire signed [DEBIT:0] score_3_x67;
wire signed [DEBIT:0] score_3_x68;
wire signed [DEBIT:0] score_3_x69;
wire signed [DEBIT:0] score_3_x70;
wire signed [DEBIT:0] score_3_x71;
wire signed [DEBIT:0] score_3_x72;
wire signed [DEBIT:0] score_3_x73;
wire signed [DEBIT:0] score_3_x74;
wire signed [DEBIT:0] score_3_x75;
wire signed [DEBIT:0] score_3_x76;
wire signed [DEBIT:0] score_3_x77;
wire signed [DEBIT:0] score_3_x78;
wire signed [DEBIT:0] score_3_x79;
wire signed [DEBIT:0] score_3_x80;
wire signed [DEBIT:0] score_3_x81;
wire signed [DEBIT:0] score_3_x82;
wire signed [DEBIT:0] score_3_x83;
wire signed [DEBIT:0] score_3_x84;
wire signed [DEBIT:0] score_3_x85;
wire signed [DEBIT:0] score_3_x86;
wire signed [DEBIT:0] score_3_x87;
wire signed [DEBIT:0] score_3_x88;
wire signed [DEBIT:0] score_3_x89;
wire signed [DEBIT:0] score_3_x90;
wire signed [DEBIT:0] score_3_x91;
wire signed [DEBIT:0] score_3_x92;
wire signed [DEBIT:0] score_3_x93;
wire signed [DEBIT:0] score_3_x94;
wire signed [DEBIT:0] score_3_x95;
wire signed [DEBIT:0] score_3_x96;
wire signed [DEBIT:0] score_3_x97;
wire signed [DEBIT:0] score_3_x98;
wire signed [DEBIT:0] score_3_x99;
wire signed [DEBIT:0] score_3_x100;
wire signed [DEBIT:0] score_3_x101;
wire signed [DEBIT:0] score_3_x102;
wire signed [DEBIT:0] score_3_x103;
wire signed [DEBIT:0] score_3_x104;
wire signed [DEBIT:0] score_3_x105;
wire signed [DEBIT:0] score_3_x106;
wire signed [DEBIT:0] score_3_x107;
wire signed [DEBIT:0] score_3_x108;
wire signed [DEBIT:0] score_3_x109;
wire signed [DEBIT:0] score_3_x110;
wire signed [DEBIT:0] score_3_x111;
wire signed [DEBIT:0] score_3_x112;
wire signed [DEBIT:0] score_3_x113;
wire signed [DEBIT:0] score_3_x114;
wire signed [DEBIT:0] score_3_x115;
wire signed [DEBIT:0] score_3_x116;
wire signed [DEBIT:0] score_3_x117;
wire signed [DEBIT:0] score_3_x118;
wire signed [DEBIT:0] score_3_x119;
wire signed [DEBIT:0] score_3_x120;
wire signed [DEBIT:0] score_3_x121;
wire signed [DEBIT:0] score_3_x122;
wire signed [DEBIT:0] score_3_x123;
wire signed [DEBIT:0] score_3_x124;
wire signed [DEBIT:0] score_3_x125;
wire signed [DEBIT:0] score_3_x126;
wire signed [DEBIT:0] score_3_x127;
wire signed [DEBIT:0] score_3_x128;
wire signed [DEBIT:0] score_3_x129;
wire signed [DEBIT:0] score_3_x130;
wire signed [DEBIT:0] score_3_x131;
wire signed [DEBIT:0] score_3_x132;
wire signed [DEBIT:0] score_3_x133;
wire signed [DEBIT:0] score_3_x134;
wire signed [DEBIT:0] score_3_x135;
wire signed [DEBIT:0] score_3_x136;
wire signed [DEBIT:0] score_3_x137;
wire signed [DEBIT:0] score_3_x138;
wire signed [DEBIT:0] score_3_x139;
wire signed [DEBIT:0] score_3_x140;
wire signed [DEBIT:0] score_3_x141;
wire signed [DEBIT:0] score_3_x142;
wire signed [DEBIT:0] score_3_x143;
wire signed [DEBIT:0] score_3_x144;
wire signed [DEBIT:0] score_3_x145;
wire signed [DEBIT:0] score_3_x146;
wire signed [DEBIT:0] score_3_x147;
wire signed [DEBIT:0] score_3_x148;
wire signed [DEBIT:0] score_3_x149;
wire signed [DEBIT:0] score_3_x150;
wire signed [DEBIT:0] score_3_x151;
wire signed [DEBIT:0] score_3_x152;
wire signed [DEBIT:0] score_3_x153;
wire signed [DEBIT:0] score_3_x154;
wire signed [DEBIT:0] score_3_x155;
wire signed [DEBIT:0] score_3_x156;
wire signed [DEBIT:0] score_3_x157;
wire signed [DEBIT:0] score_3_x158;
wire signed [DEBIT:0] score_3_x159;
wire signed [DEBIT:0] score_3_x160;
wire signed [DEBIT:0] score_3_x161;
wire signed [DEBIT:0] score_3_x162;
wire signed [DEBIT:0] score_3_x163;
wire signed [DEBIT:0] score_3_x164;
wire signed [DEBIT:0] score_3_x165;
wire signed [DEBIT:0] score_3_x166;
wire signed [DEBIT:0] score_3_x167;
wire signed [DEBIT:0] score_3_x168;
wire signed [DEBIT:0] score_3_x169;
wire signed [DEBIT:0] score_3_x170;
wire signed [DEBIT:0] score_3_x171;
wire signed [DEBIT:0] score_3_x172;
wire signed [DEBIT:0] score_3_x173;
wire signed [DEBIT:0] score_3_x174;
wire signed [DEBIT:0] score_3_x175;
wire signed [DEBIT:0] score_3_x176;
wire signed [DEBIT:0] score_3_x177;
wire signed [DEBIT:0] score_3_x178;
wire signed [DEBIT:0] score_3_x179;
wire signed [DEBIT:0] score_3_x180;
wire signed [DEBIT:0] score_3_x181;
wire signed [DEBIT:0] score_3_x182;
wire signed [DEBIT:0] score_3_x183;
wire signed [DEBIT:0] score_3_x184;
wire signed [DEBIT:0] score_3_x185;
wire signed [DEBIT:0] score_3_x186;
wire signed [DEBIT:0] score_3_x187;
wire signed [DEBIT:0] score_3_x188;
wire signed [DEBIT:0] score_3_x189;
wire signed [DEBIT:0] score_3_x190;
wire signed [DEBIT:0] score_3_x191;
wire signed [DEBIT:0] score_3_x192;
wire signed [DEBIT:0] score_3_x193;
wire signed [DEBIT:0] score_3_x194;
wire signed [DEBIT:0] score_3_x195;
wire signed [DEBIT:0] score_3_x196;
wire signed [DEBIT:0] score_3_x197;
wire signed [DEBIT:0] score_3_x198;
wire signed [DEBIT:0] score_3_x199;
wire signed [DEBIT:0] score_3_x200;
wire signed [DEBIT:0] score_3_x201;
wire signed [DEBIT:0] score_3_x202;
wire signed [DEBIT:0] score_3_x203;
wire signed [DEBIT:0] score_3_x204;
wire signed [DEBIT:0] score_3_x205;
wire signed [DEBIT:0] score_3_x206;
wire signed [DEBIT:0] score_3_x207;
wire signed [DEBIT:0] score_3_x208;
wire signed [DEBIT:0] score_3_x209;
wire signed [DEBIT:0] score_3_x210;
wire signed [DEBIT:0] score_3_x211;
wire signed [DEBIT:0] score_3_x212;
wire signed [DEBIT:0] score_3_x213;
wire signed [DEBIT:0] score_3_x214;
wire signed [DEBIT:0] score_3_x215;
wire signed [DEBIT:0] score_3_x216;
wire signed [DEBIT:0] score_3_x217;
wire signed [DEBIT:0] score_3_x218;
wire signed [DEBIT:0] score_3_x219;
wire signed [DEBIT:0] score_3_x220;
wire signed [DEBIT:0] score_3_x221;
wire signed [DEBIT:0] score_3_x222;
wire signed [DEBIT:0] score_3_x223;
wire signed [DEBIT:0] score_3_x224;
wire signed [DEBIT:0] score_3_x225;
wire signed [DEBIT:0] score_3_x226;
wire signed [DEBIT:0] score_3_x227;
wire signed [DEBIT:0] score_3_x228;
wire signed [DEBIT:0] score_3_x229;
wire signed [DEBIT:0] score_3_x230;
wire signed [DEBIT:0] score_3_x231;
wire signed [DEBIT:0] score_3_x232;
wire signed [DEBIT:0] score_3_x233;
wire signed [DEBIT:0] score_3_x234;
wire signed [DEBIT:0] score_3_x235;
wire signed [DEBIT:0] score_3_x236;
wire signed [DEBIT:0] score_3_x237;
wire signed [DEBIT:0] score_3_x238;
wire signed [DEBIT:0] score_3_x239;
wire signed [DEBIT:0] score_3_x240;
wire signed [DEBIT:0] score_3_x241;
wire signed [DEBIT:0] score_3_x242;
wire signed [DEBIT:0] score_3_x243;
wire signed [DEBIT:0] score_3_x244;
wire signed [DEBIT:0] score_3_x245;
wire signed [DEBIT:0] score_3_x246;
wire signed [DEBIT:0] score_3_x247;
wire signed [DEBIT:0] score_3_x248;
wire signed [DEBIT:0] score_3_x249;
wire signed [DEBIT:0] score_3_x250;
wire signed [DEBIT:0] score_3_x251;
wire signed [DEBIT:0] score_3_x252;
wire signed [DEBIT:0] score_3_x253;
wire signed [DEBIT:0] score_3_x254;
wire signed [DEBIT:0] score_3_x255;
wire signed [DEBIT:0] score_3_x256;
wire signed [DEBIT:0] score_3_x257;
wire signed [DEBIT:0] score_3_x258;
wire signed [DEBIT:0] score_3_x259;
wire signed [DEBIT:0] score_3_x260;
wire signed [DEBIT:0] score_3_x261;
wire signed [DEBIT:0] score_3_x262;
wire signed [DEBIT:0] score_3_x263;
wire signed [DEBIT:0] score_3_x264;
wire signed [DEBIT:0] score_3_x265;
wire signed [DEBIT:0] score_3_x266;
wire signed [DEBIT:0] score_3_x267;
wire signed [DEBIT:0] score_3_x268;
wire signed [DEBIT:0] score_3_x269;
wire signed [DEBIT:0] score_3_x270;
wire signed [DEBIT:0] score_3_x271;
wire signed [DEBIT:0] score_3_x272;
wire signed [DEBIT:0] score_3_x273;
wire signed [DEBIT:0] score_3_x274;
wire signed [DEBIT:0] score_3_x275;
wire signed [DEBIT:0] score_3_x276;
wire signed [DEBIT:0] score_3_x277;
wire signed [DEBIT:0] score_3_x278;
wire signed [DEBIT:0] score_3_x279;
wire signed [DEBIT:0] score_3_x280;
wire signed [DEBIT:0] score_3_x281;
wire signed [DEBIT:0] score_3_x282;
wire signed [DEBIT:0] score_3_x283;
wire signed [DEBIT:0] score_3_x284;
wire signed [DEBIT:0] score_3_x285;
wire signed [DEBIT:0] score_3_x286;
wire signed [DEBIT:0] score_3_x287;
wire signed [DEBIT:0] score_3_x288;
wire signed [DEBIT:0] score_3_x289;
wire signed [DEBIT:0] score_3_x290;
wire signed [DEBIT:0] score_3_x291;
wire signed [DEBIT:0] score_3_x292;
wire signed [DEBIT:0] score_3_x293;
wire signed [DEBIT:0] score_3_x294;
wire signed [DEBIT:0] score_3_x295;
wire signed [DEBIT:0] score_3_x296;
wire signed [DEBIT:0] score_3_x297;
wire signed [DEBIT:0] score_3_x298;
wire signed [DEBIT:0] score_3_x299;
wire signed [DEBIT:0] score_3_x300;
wire signed [DEBIT:0] score_3_x301;
wire signed [DEBIT:0] score_3_x302;
wire signed [DEBIT:0] score_3_x303;
wire signed [DEBIT:0] score_3_x304;
wire signed [DEBIT:0] score_3_x305;
wire signed [DEBIT:0] score_3_x306;
wire signed [DEBIT:0] score_3_x307;
wire signed [DEBIT:0] score_3_x308;
wire signed [DEBIT:0] score_3_x309;
wire signed [DEBIT:0] score_3_x310;
wire signed [DEBIT:0] score_3_x311;
wire signed [DEBIT:0] score_3_x312;
wire signed [DEBIT:0] score_3_x313;
wire signed [DEBIT:0] score_3_x314;
wire signed [DEBIT:0] score_3_x315;
wire signed [DEBIT:0] score_3_x316;
wire signed [DEBIT:0] score_3_x317;
wire signed [DEBIT:0] score_3_x318;
wire signed [DEBIT:0] score_3_x319;
wire signed [DEBIT:0] score_3_x320;
wire signed [DEBIT:0] score_3_x321;
wire signed [DEBIT:0] score_3_x322;
wire signed [DEBIT:0] score_3_x323;
wire signed [DEBIT:0] score_3_x324;
wire signed [DEBIT:0] score_3_x325;
wire signed [DEBIT:0] score_3_x326;
wire signed [DEBIT:0] score_3_x327;
wire signed [DEBIT:0] score_3_x328;
wire signed [DEBIT:0] score_3_x329;
wire signed [DEBIT:0] score_3_x330;
wire signed [DEBIT:0] score_3_x331;
wire signed [DEBIT:0] score_3_x332;
wire signed [DEBIT:0] score_3_x333;
wire signed [DEBIT:0] score_3_x334;
wire signed [DEBIT:0] score_3_x335;
wire signed [DEBIT:0] score_3_x336;
wire signed [DEBIT:0] score_3_x337;
wire signed [DEBIT:0] score_3_x338;
wire signed [DEBIT:0] score_3_x339;
wire signed [DEBIT:0] score_3_x340;
wire signed [DEBIT:0] score_3_x341;
wire signed [DEBIT:0] score_3_x342;
wire signed [DEBIT:0] score_3_x343;
wire signed [DEBIT:0] score_3_x344;
wire signed [DEBIT:0] score_3_x345;
wire signed [DEBIT:0] score_3_x346;
wire signed [DEBIT:0] score_3_x347;
wire signed [DEBIT:0] score_3_x348;
wire signed [DEBIT:0] score_3_x349;
wire signed [DEBIT:0] score_3_x350;
wire signed [DEBIT:0] score_3_x351;
wire signed [DEBIT:0] score_3_x352;
wire signed [DEBIT:0] score_3_x353;
wire signed [DEBIT:0] score_3_x354;
wire signed [DEBIT:0] score_3_x355;
wire signed [DEBIT:0] score_3_x356;
wire signed [DEBIT:0] score_3_x357;
wire signed [DEBIT:0] score_3_x358;
wire signed [DEBIT:0] score_3_x359;
wire signed [DEBIT:0] score_3_x360;
wire signed [DEBIT:0] score_3_x361;
wire signed [DEBIT:0] score_3_x362;
wire signed [DEBIT:0] score_3_x363;
wire signed [DEBIT:0] score_3_x364;
wire signed [DEBIT:0] score_3_x365;
wire signed [DEBIT:0] score_3_x366;
wire signed [DEBIT:0] score_3_x367;
wire signed [DEBIT:0] score_3_x368;
wire signed [DEBIT:0] score_3_x369;
wire signed [DEBIT:0] score_3_x370;
wire signed [DEBIT:0] score_3_x371;
wire signed [DEBIT:0] score_3_x372;
wire signed [DEBIT:0] score_3_x373;
wire signed [DEBIT:0] score_3_x374;
wire signed [DEBIT:0] score_3_x375;
wire signed [DEBIT:0] score_3_x376;
wire signed [DEBIT:0] score_3_x377;
wire signed [DEBIT:0] score_3_x378;
wire signed [DEBIT:0] score_3_x379;
wire signed [DEBIT:0] score_3_x380;
wire signed [DEBIT:0] score_3_x381;
wire signed [DEBIT:0] score_3_x382;
wire signed [DEBIT:0] score_3_x383;
wire signed [DEBIT:0] score_3_x384;
wire signed [DEBIT:0] score_3_x385;
wire signed [DEBIT:0] score_3_x386;
wire signed [DEBIT:0] score_3_x387;
wire signed [DEBIT:0] score_3_x388;
wire signed [DEBIT:0] score_3_x389;
wire signed [DEBIT:0] score_3_x390;
wire signed [DEBIT:0] score_3_x391;
wire signed [DEBIT:0] score_3_x392;
wire signed [DEBIT:0] score_3_x393;
wire signed [DEBIT:0] score_3_x394;
wire signed [DEBIT:0] score_3_x395;
wire signed [DEBIT:0] score_3_x396;
wire signed [DEBIT:0] score_3_x397;
wire signed [DEBIT:0] score_3_x398;
wire signed [DEBIT:0] score_3_x399;
wire signed [DEBIT:0] score_3_x400;
wire signed [DEBIT:0] score_3_x401;
wire signed [DEBIT:0] score_3_x402;
wire signed [DEBIT:0] score_3_x403;
wire signed [DEBIT:0] score_3_x404;
wire signed [DEBIT:0] score_3_x405;
wire signed [DEBIT:0] score_3_x406;
wire signed [DEBIT:0] score_3_x407;
wire signed [DEBIT:0] score_3_x408;
wire signed [DEBIT:0] score_3_x409;
wire signed [DEBIT:0] score_3_x410;
wire signed [DEBIT:0] score_3_x411;
wire signed [DEBIT:0] score_3_x412;
wire signed [DEBIT:0] score_3_x413;
wire signed [DEBIT:0] score_3_x414;
wire signed [DEBIT:0] score_3_x415;
wire signed [DEBIT:0] score_3_x416;
wire signed [DEBIT:0] score_3_x417;
wire signed [DEBIT:0] score_3_x418;
wire signed [DEBIT:0] score_3_x419;
wire signed [DEBIT:0] score_3_x420;
wire signed [DEBIT:0] score_3_x421;
wire signed [DEBIT:0] score_3_x422;
wire signed [DEBIT:0] score_3_x423;
wire signed [DEBIT:0] score_3_x424;
wire signed [DEBIT:0] score_3_x425;
wire signed [DEBIT:0] score_3_x426;
wire signed [DEBIT:0] score_3_x427;
wire signed [DEBIT:0] score_3_x428;
wire signed [DEBIT:0] score_3_x429;
wire signed [DEBIT:0] score_3_x430;
wire signed [DEBIT:0] score_3_x431;
wire signed [DEBIT:0] score_3_x432;
wire signed [DEBIT:0] score_3_x433;
wire signed [DEBIT:0] score_3_x434;
wire signed [DEBIT:0] score_3_x435;
wire signed [DEBIT:0] score_3_x436;
wire signed [DEBIT:0] score_3_x437;
wire signed [DEBIT:0] score_3_x438;
wire signed [DEBIT:0] score_3_x439;
wire signed [DEBIT:0] score_3_x440;
wire signed [DEBIT:0] score_3_x441;
wire signed [DEBIT:0] score_3_x442;
wire signed [DEBIT:0] score_3_x443;
wire signed [DEBIT:0] score_3_x444;
wire signed [DEBIT:0] score_3_x445;
wire signed [DEBIT:0] score_3_x446;
wire signed [DEBIT:0] score_3_x447;
wire signed [DEBIT:0] score_3_x448;
wire signed [DEBIT:0] score_3_x449;
wire signed [DEBIT:0] score_3_x450;
wire signed [DEBIT:0] score_3_x451;
wire signed [DEBIT:0] score_3_x452;
wire signed [DEBIT:0] score_3_x453;
wire signed [DEBIT:0] score_3_x454;
wire signed [DEBIT:0] score_3_x455;
wire signed [DEBIT:0] score_3_x456;
wire signed [DEBIT:0] score_3_x457;
wire signed [DEBIT:0] score_3_x458;
wire signed [DEBIT:0] score_3_x459;
wire signed [DEBIT:0] score_3_x460;
wire signed [DEBIT:0] score_3_x461;
wire signed [DEBIT:0] score_3_x462;
wire signed [DEBIT:0] score_3_x463;
wire signed [DEBIT:0] score_3_x464;
wire signed [DEBIT:0] score_3_x465;
wire signed [DEBIT:0] score_3_x466;
wire signed [DEBIT:0] score_3_x467;
wire signed [DEBIT:0] score_3_x468;
wire signed [DEBIT:0] score_3_x469;
wire signed [DEBIT:0] score_3_x470;
wire signed [DEBIT:0] score_3_x471;
wire signed [DEBIT:0] score_3_x472;
wire signed [DEBIT:0] score_3_x473;
wire signed [DEBIT:0] score_3_x474;
wire signed [DEBIT:0] score_3_x475;
wire signed [DEBIT:0] score_3_x476;
wire signed [DEBIT:0] score_3_x477;
wire signed [DEBIT:0] score_3_x478;
wire signed [DEBIT:0] score_3_x479;
wire signed [DEBIT:0] score_3_x480;
wire signed [DEBIT:0] score_3_x481;
wire signed [DEBIT:0] score_3_x482;
wire signed [DEBIT:0] score_3_x483;
wire signed [DEBIT:0] score_3_x484;
wire signed [DEBIT:0] score_3_x485;
wire signed [DEBIT:0] score_3_x486;
wire signed [DEBIT:0] score_3_x487;
wire signed [DEBIT:0] score_3_x488;
wire signed [DEBIT:0] score_3_x489;
wire signed [DEBIT:0] score_3_x490;
wire signed [DEBIT:0] score_3_x491;
wire signed [DEBIT:0] score_3_x492;
wire signed [DEBIT:0] score_3_x493;
wire signed [DEBIT:0] score_3_x494;
wire signed [DEBIT:0] score_3_x495;
wire signed [DEBIT:0] score_3_x496;
wire signed [DEBIT:0] score_3_x497;
wire signed [DEBIT:0] score_3_x498;
wire signed [DEBIT:0] score_3_x499;
wire signed [DEBIT:0] score_3_x500;
wire signed [DEBIT:0] score_3_x501;
wire signed [DEBIT:0] score_3_x502;
wire signed [DEBIT:0] score_3_x503;
wire signed [DEBIT:0] score_3_x504;
wire signed [DEBIT:0] score_3_x505;
wire signed [DEBIT:0] score_3_x506;
wire signed [DEBIT:0] score_3_x507;
wire signed [DEBIT:0] score_3_x508;
wire signed [DEBIT:0] score_3_x509;
wire signed [DEBIT:0] score_3_x510;
wire signed [DEBIT:0] score_3_x511;
wire signed [DEBIT:0] score_3_x512;
wire signed [DEBIT:0] score_3_x513;
wire signed [DEBIT:0] score_3_x514;
wire signed [DEBIT:0] score_3_x515;
wire signed [DEBIT:0] score_3_x516;
wire signed [DEBIT:0] score_3_x517;
wire signed [DEBIT:0] score_3_x518;
wire signed [DEBIT:0] score_3_x519;
wire signed [DEBIT:0] score_3_x520;
wire signed [DEBIT:0] score_3_x521;
wire signed [DEBIT:0] score_3_x522;
wire signed [DEBIT:0] score_3_x523;
wire signed [DEBIT:0] score_3_x524;
wire signed [DEBIT:0] score_3_x525;
wire signed [DEBIT:0] score_3_x526;
wire signed [DEBIT:0] score_3_x527;
wire signed [DEBIT:0] score_3_x528;
wire signed [DEBIT:0] score_3_x529;
wire signed [DEBIT:0] score_3_x530;
wire signed [DEBIT:0] score_3_x531;
wire signed [DEBIT:0] score_3_x532;
wire signed [DEBIT:0] score_3_x533;
wire signed [DEBIT:0] score_3_x534;
wire signed [DEBIT:0] score_3_x535;
wire signed [DEBIT:0] score_3_x536;
wire signed [DEBIT:0] score_3_x537;
wire signed [DEBIT:0] score_3_x538;
wire signed [DEBIT:0] score_3_x539;
wire signed [DEBIT:0] score_3_x540;
wire signed [DEBIT:0] score_3_x541;
wire signed [DEBIT:0] score_3_x542;
wire signed [DEBIT:0] score_3_x543;
wire signed [DEBIT:0] score_3_x544;
wire signed [DEBIT:0] score_3_x545;
wire signed [DEBIT:0] score_3_x546;
wire signed [DEBIT:0] score_3_x547;
wire signed [DEBIT:0] score_3_x548;
wire signed [DEBIT:0] score_3_x549;
wire signed [DEBIT:0] score_3_x550;
wire signed [DEBIT:0] score_3_x551;
wire signed [DEBIT:0] score_3_x552;
wire signed [DEBIT:0] score_3_x553;
wire signed [DEBIT:0] score_3_x554;
wire signed [DEBIT:0] score_3_x555;
wire signed [DEBIT:0] score_3_x556;
wire signed [DEBIT:0] score_3_x557;
wire signed [DEBIT:0] score_3_x558;
wire signed [DEBIT:0] score_3_x559;
wire signed [DEBIT:0] score_3_x560;
wire signed [DEBIT:0] score_3_x561;
wire signed [DEBIT:0] score_3_x562;
wire signed [DEBIT:0] score_3_x563;
wire signed [DEBIT:0] score_3_x564;
wire signed [DEBIT:0] score_3_x565;
wire signed [DEBIT:0] score_3_x566;
wire signed [DEBIT:0] score_3_x567;
wire signed [DEBIT:0] score_3_x568;
wire signed [DEBIT:0] score_3_x569;
wire signed [DEBIT:0] score_3_x570;
wire signed [DEBIT:0] score_3_x571;
wire signed [DEBIT:0] score_3_x572;
wire signed [DEBIT:0] score_3_x573;
wire signed [DEBIT:0] score_3_x574;
wire signed [DEBIT:0] score_3_x575;
wire signed [DEBIT:0] score_3_x576;
wire signed [DEBIT:0] score_3_x577;
wire signed [DEBIT:0] score_3_x578;
wire signed [DEBIT:0] score_3_x579;
wire signed [DEBIT:0] score_3_x580;
wire signed [DEBIT:0] score_3_x581;
wire signed [DEBIT:0] score_3_x582;
wire signed [DEBIT:0] score_3_x583;
wire signed [DEBIT:0] score_3_x584;
wire signed [DEBIT:0] score_3_x585;
wire signed [DEBIT:0] score_3_x586;
wire signed [DEBIT:0] score_3_x587;
wire signed [DEBIT:0] score_3_x588;
wire signed [DEBIT:0] score_3_x589;
wire signed [DEBIT:0] score_3_x590;
wire signed [DEBIT:0] score_3_x591;
wire signed [DEBIT:0] score_3_x592;
wire signed [DEBIT:0] score_3_x593;
wire signed [DEBIT:0] score_3_x594;
wire signed [DEBIT:0] score_3_x595;
wire signed [DEBIT:0] score_3_x596;
wire signed [DEBIT:0] score_3_x597;
wire signed [DEBIT:0] score_3_x598;
wire signed [DEBIT:0] score_3_x599;
wire signed [DEBIT:0] score_3_x600;
wire signed [DEBIT:0] score_3_x601;
wire signed [DEBIT:0] score_3_x602;
wire signed [DEBIT:0] score_3_x603;
wire signed [DEBIT:0] score_3_x604;
wire signed [DEBIT:0] score_3_x605;
wire signed [DEBIT:0] score_3_x606;
wire signed [DEBIT:0] score_3_x607;
wire signed [DEBIT:0] score_3_x608;
wire signed [DEBIT:0] score_3_x609;
wire signed [DEBIT:0] score_3_x610;
wire signed [DEBIT:0] score_3_x611;
wire signed [DEBIT:0] score_3_x612;
wire signed [DEBIT:0] score_3_x613;
wire signed [DEBIT:0] score_3_x614;
wire signed [DEBIT:0] score_3_x615;
wire signed [DEBIT:0] score_3_x616;
wire signed [DEBIT:0] score_3_x617;
wire signed [DEBIT:0] score_3_x618;
wire signed [DEBIT:0] score_3_x619;
wire signed [DEBIT:0] score_3_x620;
wire signed [DEBIT:0] score_3_x621;
wire signed [DEBIT:0] score_3_x622;
wire signed [DEBIT:0] score_3_x623;
wire signed [DEBIT:0] score_3_x624;
wire signed [DEBIT:0] score_3_x625;
wire signed [DEBIT:0] score_3_x626;
wire signed [DEBIT:0] score_3_x627;
wire signed [DEBIT:0] score_3_x628;
wire signed [DEBIT:0] score_3_x629;
wire signed [DEBIT:0] score_3_x630;
wire signed [DEBIT:0] score_3_x631;
wire signed [DEBIT:0] score_3_x632;
wire signed [DEBIT:0] score_3_x633;
wire signed [DEBIT:0] score_3_x634;
wire signed [DEBIT:0] score_3_x635;
wire signed [DEBIT:0] score_3_x636;
wire signed [DEBIT:0] score_3_x637;
wire signed [DEBIT:0] score_3_x638;
wire signed [DEBIT:0] score_3_x639;
wire signed [DEBIT:0] score_3_x640;
wire signed [DEBIT:0] score_3_x641;
wire signed [DEBIT:0] score_3_x642;
wire signed [DEBIT:0] score_3_x643;
wire signed [DEBIT:0] score_3_x644;
wire signed [DEBIT:0] score_3_x645;
wire signed [DEBIT:0] score_3_x646;
wire signed [DEBIT:0] score_3_x647;
wire signed [DEBIT:0] score_3_x648;
wire signed [DEBIT:0] score_3_x649;
wire signed [DEBIT:0] score_3_x650;
wire signed [DEBIT:0] score_3_x651;
wire signed [DEBIT:0] score_3_x652;
wire signed [DEBIT:0] score_3_x653;
wire signed [DEBIT:0] score_3_x654;
wire signed [DEBIT:0] score_3_x655;
wire signed [DEBIT:0] score_3_x656;
wire signed [DEBIT:0] score_3_x657;
wire signed [DEBIT:0] score_3_x658;
wire signed [DEBIT:0] score_3_x659;
wire signed [DEBIT:0] score_3_x660;
wire signed [DEBIT:0] score_3_x661;
wire signed [DEBIT:0] score_3_x662;
wire signed [DEBIT:0] score_3_x663;
wire signed [DEBIT:0] score_3_x664;
wire signed [DEBIT:0] score_3_x665;
wire signed [DEBIT:0] score_3_x666;
wire signed [DEBIT:0] score_3_x667;
wire signed [DEBIT:0] score_3_x668;
wire signed [DEBIT:0] score_3_x669;
wire signed [DEBIT:0] score_3_x670;
wire signed [DEBIT:0] score_3_x671;
wire signed [DEBIT:0] score_3_x672;
wire signed [DEBIT:0] score_3_x673;
wire signed [DEBIT:0] score_3_x674;
wire signed [DEBIT:0] score_3_x675;
wire signed [DEBIT:0] score_3_x676;
wire signed [DEBIT:0] score_3_x677;
wire signed [DEBIT:0] score_3_x678;
wire signed [DEBIT:0] score_3_x679;
wire signed [DEBIT:0] score_3_x680;
wire signed [DEBIT:0] score_3_x681;
wire signed [DEBIT:0] score_3_x682;
wire signed [DEBIT:0] score_3_x683;
wire signed [DEBIT:0] score_3_x684;
wire signed [DEBIT:0] score_3_x685;
wire signed [DEBIT:0] score_3_x686;
wire signed [DEBIT:0] score_3_x687;
wire signed [DEBIT:0] score_3_x688;
wire signed [DEBIT:0] score_3_x689;
wire signed [DEBIT:0] score_3_x690;
wire signed [DEBIT:0] score_3_x691;
wire signed [DEBIT:0] score_3_x692;
wire signed [DEBIT:0] score_3_x693;
wire signed [DEBIT:0] score_3_x694;
wire signed [DEBIT:0] score_3_x695;
wire signed [DEBIT:0] score_3_x696;
wire signed [DEBIT:0] score_3_x697;
wire signed [DEBIT:0] score_3_x698;
wire signed [DEBIT:0] score_3_x699;
wire signed [DEBIT:0] score_3_x700;
wire signed [DEBIT:0] score_3_x701;
wire signed [DEBIT:0] score_3_x702;
wire signed [DEBIT:0] score_3_x703;
wire signed [DEBIT:0] score_3_x704;
wire signed [DEBIT:0] score_3_x705;
wire signed [DEBIT:0] score_3_x706;
wire signed [DEBIT:0] score_3_x707;
wire signed [DEBIT:0] score_3_x708;
wire signed [DEBIT:0] score_3_x709;
wire signed [DEBIT:0] score_3_x710;
wire signed [DEBIT:0] score_3_x711;
wire signed [DEBIT:0] score_3_x712;
wire signed [DEBIT:0] score_3_x713;
wire signed [DEBIT:0] score_3_x714;
wire signed [DEBIT:0] score_3_x715;
wire signed [DEBIT:0] score_3_x716;
wire signed [DEBIT:0] score_3_x717;
wire signed [DEBIT:0] score_3_x718;
wire signed [DEBIT:0] score_3_x719;
wire signed [DEBIT:0] score_3_x720;
wire signed [DEBIT:0] score_3_x721;
wire signed [DEBIT:0] score_3_x722;
wire signed [DEBIT:0] score_3_x723;
wire signed [DEBIT:0] score_3_x724;
wire signed [DEBIT:0] score_3_x725;
wire signed [DEBIT:0] score_3_x726;
wire signed [DEBIT:0] score_3_x727;
wire signed [DEBIT:0] score_3_x728;
wire signed [DEBIT:0] score_3_x729;
wire signed [DEBIT:0] score_3_x730;
wire signed [DEBIT:0] score_3_x731;
wire signed [DEBIT:0] score_3_x732;
wire signed [DEBIT:0] score_3_x733;
wire signed [DEBIT:0] score_3_x734;
wire signed [DEBIT:0] score_3_x735;
wire signed [DEBIT:0] score_3_x736;
wire signed [DEBIT:0] score_3_x737;
wire signed [DEBIT:0] score_3_x738;
wire signed [DEBIT:0] score_3_x739;
wire signed [DEBIT:0] score_3_x740;
wire signed [DEBIT:0] score_3_x741;
wire signed [DEBIT:0] score_3_x742;
wire signed [DEBIT:0] score_3_x743;
wire signed [DEBIT:0] score_3_x744;
wire signed [DEBIT:0] score_3_x745;
wire signed [DEBIT:0] score_3_x746;
wire signed [DEBIT:0] score_3_x747;
wire signed [DEBIT:0] score_3_x748;
wire signed [DEBIT:0] score_3_x749;
wire signed [DEBIT:0] score_3_x750;
wire signed [DEBIT:0] score_3_x751;
wire signed [DEBIT:0] score_3_x752;
wire signed [DEBIT:0] score_3_x753;
wire signed [DEBIT:0] score_3_x754;
wire signed [DEBIT:0] score_3_x755;
wire signed [DEBIT:0] score_3_x756;
wire signed [DEBIT:0] score_3_x757;
wire signed [DEBIT:0] score_3_x758;
wire signed [DEBIT:0] score_3_x759;
wire signed [DEBIT:0] score_3_x760;
wire signed [DEBIT:0] score_3_x761;
wire signed [DEBIT:0] score_3_x762;
wire signed [DEBIT:0] score_3_x763;
wire signed [DEBIT:0] score_3_x764;
wire signed [DEBIT:0] score_3_x765;
wire signed [DEBIT:0] score_3_x766;
wire signed [DEBIT:0] score_3_x767;
wire signed [DEBIT:0] score_3_x768;
wire signed [DEBIT:0] score_3_x769;
wire signed [DEBIT:0] score_3_x770;
wire signed [DEBIT:0] score_3_x771;
wire signed [DEBIT:0] score_3_x772;
wire signed [DEBIT:0] score_3_x773;
wire signed [DEBIT:0] score_3_x774;
wire signed [DEBIT:0] score_3_x775;
wire signed [DEBIT:0] score_3_x776;
wire signed [DEBIT:0] score_3_x777;
wire signed [DEBIT:0] score_3_x778;
wire signed [DEBIT:0] score_3_x779;
wire signed [DEBIT:0] score_3_x780;
wire signed [DEBIT:0] score_3_x781;
wire signed [DEBIT:0] score_3_x782;
wire signed [DEBIT:0] score_3_x783;
wire signed [DEBIT:0] score_3_x784;
wire signed [DEBIT:0] score_4_x1;
wire signed [DEBIT:0] score_4_x2;
wire signed [DEBIT:0] score_4_x3;
wire signed [DEBIT:0] score_4_x4;
wire signed [DEBIT:0] score_4_x5;
wire signed [DEBIT:0] score_4_x6;
wire signed [DEBIT:0] score_4_x7;
wire signed [DEBIT:0] score_4_x8;
wire signed [DEBIT:0] score_4_x9;
wire signed [DEBIT:0] score_4_x10;
wire signed [DEBIT:0] score_4_x11;
wire signed [DEBIT:0] score_4_x12;
wire signed [DEBIT:0] score_4_x13;
wire signed [DEBIT:0] score_4_x14;
wire signed [DEBIT:0] score_4_x15;
wire signed [DEBIT:0] score_4_x16;
wire signed [DEBIT:0] score_4_x17;
wire signed [DEBIT:0] score_4_x18;
wire signed [DEBIT:0] score_4_x19;
wire signed [DEBIT:0] score_4_x20;
wire signed [DEBIT:0] score_4_x21;
wire signed [DEBIT:0] score_4_x22;
wire signed [DEBIT:0] score_4_x23;
wire signed [DEBIT:0] score_4_x24;
wire signed [DEBIT:0] score_4_x25;
wire signed [DEBIT:0] score_4_x26;
wire signed [DEBIT:0] score_4_x27;
wire signed [DEBIT:0] score_4_x28;
wire signed [DEBIT:0] score_4_x29;
wire signed [DEBIT:0] score_4_x30;
wire signed [DEBIT:0] score_4_x31;
wire signed [DEBIT:0] score_4_x32;
wire signed [DEBIT:0] score_4_x33;
wire signed [DEBIT:0] score_4_x34;
wire signed [DEBIT:0] score_4_x35;
wire signed [DEBIT:0] score_4_x36;
wire signed [DEBIT:0] score_4_x37;
wire signed [DEBIT:0] score_4_x38;
wire signed [DEBIT:0] score_4_x39;
wire signed [DEBIT:0] score_4_x40;
wire signed [DEBIT:0] score_4_x41;
wire signed [DEBIT:0] score_4_x42;
wire signed [DEBIT:0] score_4_x43;
wire signed [DEBIT:0] score_4_x44;
wire signed [DEBIT:0] score_4_x45;
wire signed [DEBIT:0] score_4_x46;
wire signed [DEBIT:0] score_4_x47;
wire signed [DEBIT:0] score_4_x48;
wire signed [DEBIT:0] score_4_x49;
wire signed [DEBIT:0] score_4_x50;
wire signed [DEBIT:0] score_4_x51;
wire signed [DEBIT:0] score_4_x52;
wire signed [DEBIT:0] score_4_x53;
wire signed [DEBIT:0] score_4_x54;
wire signed [DEBIT:0] score_4_x55;
wire signed [DEBIT:0] score_4_x56;
wire signed [DEBIT:0] score_4_x57;
wire signed [DEBIT:0] score_4_x58;
wire signed [DEBIT:0] score_4_x59;
wire signed [DEBIT:0] score_4_x60;
wire signed [DEBIT:0] score_4_x61;
wire signed [DEBIT:0] score_4_x62;
wire signed [DEBIT:0] score_4_x63;
wire signed [DEBIT:0] score_4_x64;
wire signed [DEBIT:0] score_4_x65;
wire signed [DEBIT:0] score_4_x66;
wire signed [DEBIT:0] score_4_x67;
wire signed [DEBIT:0] score_4_x68;
wire signed [DEBIT:0] score_4_x69;
wire signed [DEBIT:0] score_4_x70;
wire signed [DEBIT:0] score_4_x71;
wire signed [DEBIT:0] score_4_x72;
wire signed [DEBIT:0] score_4_x73;
wire signed [DEBIT:0] score_4_x74;
wire signed [DEBIT:0] score_4_x75;
wire signed [DEBIT:0] score_4_x76;
wire signed [DEBIT:0] score_4_x77;
wire signed [DEBIT:0] score_4_x78;
wire signed [DEBIT:0] score_4_x79;
wire signed [DEBIT:0] score_4_x80;
wire signed [DEBIT:0] score_4_x81;
wire signed [DEBIT:0] score_4_x82;
wire signed [DEBIT:0] score_4_x83;
wire signed [DEBIT:0] score_4_x84;
wire signed [DEBIT:0] score_4_x85;
wire signed [DEBIT:0] score_4_x86;
wire signed [DEBIT:0] score_4_x87;
wire signed [DEBIT:0] score_4_x88;
wire signed [DEBIT:0] score_4_x89;
wire signed [DEBIT:0] score_4_x90;
wire signed [DEBIT:0] score_4_x91;
wire signed [DEBIT:0] score_4_x92;
wire signed [DEBIT:0] score_4_x93;
wire signed [DEBIT:0] score_4_x94;
wire signed [DEBIT:0] score_4_x95;
wire signed [DEBIT:0] score_4_x96;
wire signed [DEBIT:0] score_4_x97;
wire signed [DEBIT:0] score_4_x98;
wire signed [DEBIT:0] score_4_x99;
wire signed [DEBIT:0] score_4_x100;
wire signed [DEBIT:0] score_4_x101;
wire signed [DEBIT:0] score_4_x102;
wire signed [DEBIT:0] score_4_x103;
wire signed [DEBIT:0] score_4_x104;
wire signed [DEBIT:0] score_4_x105;
wire signed [DEBIT:0] score_4_x106;
wire signed [DEBIT:0] score_4_x107;
wire signed [DEBIT:0] score_4_x108;
wire signed [DEBIT:0] score_4_x109;
wire signed [DEBIT:0] score_4_x110;
wire signed [DEBIT:0] score_4_x111;
wire signed [DEBIT:0] score_4_x112;
wire signed [DEBIT:0] score_4_x113;
wire signed [DEBIT:0] score_4_x114;
wire signed [DEBIT:0] score_4_x115;
wire signed [DEBIT:0] score_4_x116;
wire signed [DEBIT:0] score_4_x117;
wire signed [DEBIT:0] score_4_x118;
wire signed [DEBIT:0] score_4_x119;
wire signed [DEBIT:0] score_4_x120;
wire signed [DEBIT:0] score_4_x121;
wire signed [DEBIT:0] score_4_x122;
wire signed [DEBIT:0] score_4_x123;
wire signed [DEBIT:0] score_4_x124;
wire signed [DEBIT:0] score_4_x125;
wire signed [DEBIT:0] score_4_x126;
wire signed [DEBIT:0] score_4_x127;
wire signed [DEBIT:0] score_4_x128;
wire signed [DEBIT:0] score_4_x129;
wire signed [DEBIT:0] score_4_x130;
wire signed [DEBIT:0] score_4_x131;
wire signed [DEBIT:0] score_4_x132;
wire signed [DEBIT:0] score_4_x133;
wire signed [DEBIT:0] score_4_x134;
wire signed [DEBIT:0] score_4_x135;
wire signed [DEBIT:0] score_4_x136;
wire signed [DEBIT:0] score_4_x137;
wire signed [DEBIT:0] score_4_x138;
wire signed [DEBIT:0] score_4_x139;
wire signed [DEBIT:0] score_4_x140;
wire signed [DEBIT:0] score_4_x141;
wire signed [DEBIT:0] score_4_x142;
wire signed [DEBIT:0] score_4_x143;
wire signed [DEBIT:0] score_4_x144;
wire signed [DEBIT:0] score_4_x145;
wire signed [DEBIT:0] score_4_x146;
wire signed [DEBIT:0] score_4_x147;
wire signed [DEBIT:0] score_4_x148;
wire signed [DEBIT:0] score_4_x149;
wire signed [DEBIT:0] score_4_x150;
wire signed [DEBIT:0] score_4_x151;
wire signed [DEBIT:0] score_4_x152;
wire signed [DEBIT:0] score_4_x153;
wire signed [DEBIT:0] score_4_x154;
wire signed [DEBIT:0] score_4_x155;
wire signed [DEBIT:0] score_4_x156;
wire signed [DEBIT:0] score_4_x157;
wire signed [DEBIT:0] score_4_x158;
wire signed [DEBIT:0] score_4_x159;
wire signed [DEBIT:0] score_4_x160;
wire signed [DEBIT:0] score_4_x161;
wire signed [DEBIT:0] score_4_x162;
wire signed [DEBIT:0] score_4_x163;
wire signed [DEBIT:0] score_4_x164;
wire signed [DEBIT:0] score_4_x165;
wire signed [DEBIT:0] score_4_x166;
wire signed [DEBIT:0] score_4_x167;
wire signed [DEBIT:0] score_4_x168;
wire signed [DEBIT:0] score_4_x169;
wire signed [DEBIT:0] score_4_x170;
wire signed [DEBIT:0] score_4_x171;
wire signed [DEBIT:0] score_4_x172;
wire signed [DEBIT:0] score_4_x173;
wire signed [DEBIT:0] score_4_x174;
wire signed [DEBIT:0] score_4_x175;
wire signed [DEBIT:0] score_4_x176;
wire signed [DEBIT:0] score_4_x177;
wire signed [DEBIT:0] score_4_x178;
wire signed [DEBIT:0] score_4_x179;
wire signed [DEBIT:0] score_4_x180;
wire signed [DEBIT:0] score_4_x181;
wire signed [DEBIT:0] score_4_x182;
wire signed [DEBIT:0] score_4_x183;
wire signed [DEBIT:0] score_4_x184;
wire signed [DEBIT:0] score_4_x185;
wire signed [DEBIT:0] score_4_x186;
wire signed [DEBIT:0] score_4_x187;
wire signed [DEBIT:0] score_4_x188;
wire signed [DEBIT:0] score_4_x189;
wire signed [DEBIT:0] score_4_x190;
wire signed [DEBIT:0] score_4_x191;
wire signed [DEBIT:0] score_4_x192;
wire signed [DEBIT:0] score_4_x193;
wire signed [DEBIT:0] score_4_x194;
wire signed [DEBIT:0] score_4_x195;
wire signed [DEBIT:0] score_4_x196;
wire signed [DEBIT:0] score_4_x197;
wire signed [DEBIT:0] score_4_x198;
wire signed [DEBIT:0] score_4_x199;
wire signed [DEBIT:0] score_4_x200;
wire signed [DEBIT:0] score_4_x201;
wire signed [DEBIT:0] score_4_x202;
wire signed [DEBIT:0] score_4_x203;
wire signed [DEBIT:0] score_4_x204;
wire signed [DEBIT:0] score_4_x205;
wire signed [DEBIT:0] score_4_x206;
wire signed [DEBIT:0] score_4_x207;
wire signed [DEBIT:0] score_4_x208;
wire signed [DEBIT:0] score_4_x209;
wire signed [DEBIT:0] score_4_x210;
wire signed [DEBIT:0] score_4_x211;
wire signed [DEBIT:0] score_4_x212;
wire signed [DEBIT:0] score_4_x213;
wire signed [DEBIT:0] score_4_x214;
wire signed [DEBIT:0] score_4_x215;
wire signed [DEBIT:0] score_4_x216;
wire signed [DEBIT:0] score_4_x217;
wire signed [DEBIT:0] score_4_x218;
wire signed [DEBIT:0] score_4_x219;
wire signed [DEBIT:0] score_4_x220;
wire signed [DEBIT:0] score_4_x221;
wire signed [DEBIT:0] score_4_x222;
wire signed [DEBIT:0] score_4_x223;
wire signed [DEBIT:0] score_4_x224;
wire signed [DEBIT:0] score_4_x225;
wire signed [DEBIT:0] score_4_x226;
wire signed [DEBIT:0] score_4_x227;
wire signed [DEBIT:0] score_4_x228;
wire signed [DEBIT:0] score_4_x229;
wire signed [DEBIT:0] score_4_x230;
wire signed [DEBIT:0] score_4_x231;
wire signed [DEBIT:0] score_4_x232;
wire signed [DEBIT:0] score_4_x233;
wire signed [DEBIT:0] score_4_x234;
wire signed [DEBIT:0] score_4_x235;
wire signed [DEBIT:0] score_4_x236;
wire signed [DEBIT:0] score_4_x237;
wire signed [DEBIT:0] score_4_x238;
wire signed [DEBIT:0] score_4_x239;
wire signed [DEBIT:0] score_4_x240;
wire signed [DEBIT:0] score_4_x241;
wire signed [DEBIT:0] score_4_x242;
wire signed [DEBIT:0] score_4_x243;
wire signed [DEBIT:0] score_4_x244;
wire signed [DEBIT:0] score_4_x245;
wire signed [DEBIT:0] score_4_x246;
wire signed [DEBIT:0] score_4_x247;
wire signed [DEBIT:0] score_4_x248;
wire signed [DEBIT:0] score_4_x249;
wire signed [DEBIT:0] score_4_x250;
wire signed [DEBIT:0] score_4_x251;
wire signed [DEBIT:0] score_4_x252;
wire signed [DEBIT:0] score_4_x253;
wire signed [DEBIT:0] score_4_x254;
wire signed [DEBIT:0] score_4_x255;
wire signed [DEBIT:0] score_4_x256;
wire signed [DEBIT:0] score_4_x257;
wire signed [DEBIT:0] score_4_x258;
wire signed [DEBIT:0] score_4_x259;
wire signed [DEBIT:0] score_4_x260;
wire signed [DEBIT:0] score_4_x261;
wire signed [DEBIT:0] score_4_x262;
wire signed [DEBIT:0] score_4_x263;
wire signed [DEBIT:0] score_4_x264;
wire signed [DEBIT:0] score_4_x265;
wire signed [DEBIT:0] score_4_x266;
wire signed [DEBIT:0] score_4_x267;
wire signed [DEBIT:0] score_4_x268;
wire signed [DEBIT:0] score_4_x269;
wire signed [DEBIT:0] score_4_x270;
wire signed [DEBIT:0] score_4_x271;
wire signed [DEBIT:0] score_4_x272;
wire signed [DEBIT:0] score_4_x273;
wire signed [DEBIT:0] score_4_x274;
wire signed [DEBIT:0] score_4_x275;
wire signed [DEBIT:0] score_4_x276;
wire signed [DEBIT:0] score_4_x277;
wire signed [DEBIT:0] score_4_x278;
wire signed [DEBIT:0] score_4_x279;
wire signed [DEBIT:0] score_4_x280;
wire signed [DEBIT:0] score_4_x281;
wire signed [DEBIT:0] score_4_x282;
wire signed [DEBIT:0] score_4_x283;
wire signed [DEBIT:0] score_4_x284;
wire signed [DEBIT:0] score_4_x285;
wire signed [DEBIT:0] score_4_x286;
wire signed [DEBIT:0] score_4_x287;
wire signed [DEBIT:0] score_4_x288;
wire signed [DEBIT:0] score_4_x289;
wire signed [DEBIT:0] score_4_x290;
wire signed [DEBIT:0] score_4_x291;
wire signed [DEBIT:0] score_4_x292;
wire signed [DEBIT:0] score_4_x293;
wire signed [DEBIT:0] score_4_x294;
wire signed [DEBIT:0] score_4_x295;
wire signed [DEBIT:0] score_4_x296;
wire signed [DEBIT:0] score_4_x297;
wire signed [DEBIT:0] score_4_x298;
wire signed [DEBIT:0] score_4_x299;
wire signed [DEBIT:0] score_4_x300;
wire signed [DEBIT:0] score_4_x301;
wire signed [DEBIT:0] score_4_x302;
wire signed [DEBIT:0] score_4_x303;
wire signed [DEBIT:0] score_4_x304;
wire signed [DEBIT:0] score_4_x305;
wire signed [DEBIT:0] score_4_x306;
wire signed [DEBIT:0] score_4_x307;
wire signed [DEBIT:0] score_4_x308;
wire signed [DEBIT:0] score_4_x309;
wire signed [DEBIT:0] score_4_x310;
wire signed [DEBIT:0] score_4_x311;
wire signed [DEBIT:0] score_4_x312;
wire signed [DEBIT:0] score_4_x313;
wire signed [DEBIT:0] score_4_x314;
wire signed [DEBIT:0] score_4_x315;
wire signed [DEBIT:0] score_4_x316;
wire signed [DEBIT:0] score_4_x317;
wire signed [DEBIT:0] score_4_x318;
wire signed [DEBIT:0] score_4_x319;
wire signed [DEBIT:0] score_4_x320;
wire signed [DEBIT:0] score_4_x321;
wire signed [DEBIT:0] score_4_x322;
wire signed [DEBIT:0] score_4_x323;
wire signed [DEBIT:0] score_4_x324;
wire signed [DEBIT:0] score_4_x325;
wire signed [DEBIT:0] score_4_x326;
wire signed [DEBIT:0] score_4_x327;
wire signed [DEBIT:0] score_4_x328;
wire signed [DEBIT:0] score_4_x329;
wire signed [DEBIT:0] score_4_x330;
wire signed [DEBIT:0] score_4_x331;
wire signed [DEBIT:0] score_4_x332;
wire signed [DEBIT:0] score_4_x333;
wire signed [DEBIT:0] score_4_x334;
wire signed [DEBIT:0] score_4_x335;
wire signed [DEBIT:0] score_4_x336;
wire signed [DEBIT:0] score_4_x337;
wire signed [DEBIT:0] score_4_x338;
wire signed [DEBIT:0] score_4_x339;
wire signed [DEBIT:0] score_4_x340;
wire signed [DEBIT:0] score_4_x341;
wire signed [DEBIT:0] score_4_x342;
wire signed [DEBIT:0] score_4_x343;
wire signed [DEBIT:0] score_4_x344;
wire signed [DEBIT:0] score_4_x345;
wire signed [DEBIT:0] score_4_x346;
wire signed [DEBIT:0] score_4_x347;
wire signed [DEBIT:0] score_4_x348;
wire signed [DEBIT:0] score_4_x349;
wire signed [DEBIT:0] score_4_x350;
wire signed [DEBIT:0] score_4_x351;
wire signed [DEBIT:0] score_4_x352;
wire signed [DEBIT:0] score_4_x353;
wire signed [DEBIT:0] score_4_x354;
wire signed [DEBIT:0] score_4_x355;
wire signed [DEBIT:0] score_4_x356;
wire signed [DEBIT:0] score_4_x357;
wire signed [DEBIT:0] score_4_x358;
wire signed [DEBIT:0] score_4_x359;
wire signed [DEBIT:0] score_4_x360;
wire signed [DEBIT:0] score_4_x361;
wire signed [DEBIT:0] score_4_x362;
wire signed [DEBIT:0] score_4_x363;
wire signed [DEBIT:0] score_4_x364;
wire signed [DEBIT:0] score_4_x365;
wire signed [DEBIT:0] score_4_x366;
wire signed [DEBIT:0] score_4_x367;
wire signed [DEBIT:0] score_4_x368;
wire signed [DEBIT:0] score_4_x369;
wire signed [DEBIT:0] score_4_x370;
wire signed [DEBIT:0] score_4_x371;
wire signed [DEBIT:0] score_4_x372;
wire signed [DEBIT:0] score_4_x373;
wire signed [DEBIT:0] score_4_x374;
wire signed [DEBIT:0] score_4_x375;
wire signed [DEBIT:0] score_4_x376;
wire signed [DEBIT:0] score_4_x377;
wire signed [DEBIT:0] score_4_x378;
wire signed [DEBIT:0] score_4_x379;
wire signed [DEBIT:0] score_4_x380;
wire signed [DEBIT:0] score_4_x381;
wire signed [DEBIT:0] score_4_x382;
wire signed [DEBIT:0] score_4_x383;
wire signed [DEBIT:0] score_4_x384;
wire signed [DEBIT:0] score_4_x385;
wire signed [DEBIT:0] score_4_x386;
wire signed [DEBIT:0] score_4_x387;
wire signed [DEBIT:0] score_4_x388;
wire signed [DEBIT:0] score_4_x389;
wire signed [DEBIT:0] score_4_x390;
wire signed [DEBIT:0] score_4_x391;
wire signed [DEBIT:0] score_4_x392;
wire signed [DEBIT:0] score_4_x393;
wire signed [DEBIT:0] score_4_x394;
wire signed [DEBIT:0] score_4_x395;
wire signed [DEBIT:0] score_4_x396;
wire signed [DEBIT:0] score_4_x397;
wire signed [DEBIT:0] score_4_x398;
wire signed [DEBIT:0] score_4_x399;
wire signed [DEBIT:0] score_4_x400;
wire signed [DEBIT:0] score_4_x401;
wire signed [DEBIT:0] score_4_x402;
wire signed [DEBIT:0] score_4_x403;
wire signed [DEBIT:0] score_4_x404;
wire signed [DEBIT:0] score_4_x405;
wire signed [DEBIT:0] score_4_x406;
wire signed [DEBIT:0] score_4_x407;
wire signed [DEBIT:0] score_4_x408;
wire signed [DEBIT:0] score_4_x409;
wire signed [DEBIT:0] score_4_x410;
wire signed [DEBIT:0] score_4_x411;
wire signed [DEBIT:0] score_4_x412;
wire signed [DEBIT:0] score_4_x413;
wire signed [DEBIT:0] score_4_x414;
wire signed [DEBIT:0] score_4_x415;
wire signed [DEBIT:0] score_4_x416;
wire signed [DEBIT:0] score_4_x417;
wire signed [DEBIT:0] score_4_x418;
wire signed [DEBIT:0] score_4_x419;
wire signed [DEBIT:0] score_4_x420;
wire signed [DEBIT:0] score_4_x421;
wire signed [DEBIT:0] score_4_x422;
wire signed [DEBIT:0] score_4_x423;
wire signed [DEBIT:0] score_4_x424;
wire signed [DEBIT:0] score_4_x425;
wire signed [DEBIT:0] score_4_x426;
wire signed [DEBIT:0] score_4_x427;
wire signed [DEBIT:0] score_4_x428;
wire signed [DEBIT:0] score_4_x429;
wire signed [DEBIT:0] score_4_x430;
wire signed [DEBIT:0] score_4_x431;
wire signed [DEBIT:0] score_4_x432;
wire signed [DEBIT:0] score_4_x433;
wire signed [DEBIT:0] score_4_x434;
wire signed [DEBIT:0] score_4_x435;
wire signed [DEBIT:0] score_4_x436;
wire signed [DEBIT:0] score_4_x437;
wire signed [DEBIT:0] score_4_x438;
wire signed [DEBIT:0] score_4_x439;
wire signed [DEBIT:0] score_4_x440;
wire signed [DEBIT:0] score_4_x441;
wire signed [DEBIT:0] score_4_x442;
wire signed [DEBIT:0] score_4_x443;
wire signed [DEBIT:0] score_4_x444;
wire signed [DEBIT:0] score_4_x445;
wire signed [DEBIT:0] score_4_x446;
wire signed [DEBIT:0] score_4_x447;
wire signed [DEBIT:0] score_4_x448;
wire signed [DEBIT:0] score_4_x449;
wire signed [DEBIT:0] score_4_x450;
wire signed [DEBIT:0] score_4_x451;
wire signed [DEBIT:0] score_4_x452;
wire signed [DEBIT:0] score_4_x453;
wire signed [DEBIT:0] score_4_x454;
wire signed [DEBIT:0] score_4_x455;
wire signed [DEBIT:0] score_4_x456;
wire signed [DEBIT:0] score_4_x457;
wire signed [DEBIT:0] score_4_x458;
wire signed [DEBIT:0] score_4_x459;
wire signed [DEBIT:0] score_4_x460;
wire signed [DEBIT:0] score_4_x461;
wire signed [DEBIT:0] score_4_x462;
wire signed [DEBIT:0] score_4_x463;
wire signed [DEBIT:0] score_4_x464;
wire signed [DEBIT:0] score_4_x465;
wire signed [DEBIT:0] score_4_x466;
wire signed [DEBIT:0] score_4_x467;
wire signed [DEBIT:0] score_4_x468;
wire signed [DEBIT:0] score_4_x469;
wire signed [DEBIT:0] score_4_x470;
wire signed [DEBIT:0] score_4_x471;
wire signed [DEBIT:0] score_4_x472;
wire signed [DEBIT:0] score_4_x473;
wire signed [DEBIT:0] score_4_x474;
wire signed [DEBIT:0] score_4_x475;
wire signed [DEBIT:0] score_4_x476;
wire signed [DEBIT:0] score_4_x477;
wire signed [DEBIT:0] score_4_x478;
wire signed [DEBIT:0] score_4_x479;
wire signed [DEBIT:0] score_4_x480;
wire signed [DEBIT:0] score_4_x481;
wire signed [DEBIT:0] score_4_x482;
wire signed [DEBIT:0] score_4_x483;
wire signed [DEBIT:0] score_4_x484;
wire signed [DEBIT:0] score_4_x485;
wire signed [DEBIT:0] score_4_x486;
wire signed [DEBIT:0] score_4_x487;
wire signed [DEBIT:0] score_4_x488;
wire signed [DEBIT:0] score_4_x489;
wire signed [DEBIT:0] score_4_x490;
wire signed [DEBIT:0] score_4_x491;
wire signed [DEBIT:0] score_4_x492;
wire signed [DEBIT:0] score_4_x493;
wire signed [DEBIT:0] score_4_x494;
wire signed [DEBIT:0] score_4_x495;
wire signed [DEBIT:0] score_4_x496;
wire signed [DEBIT:0] score_4_x497;
wire signed [DEBIT:0] score_4_x498;
wire signed [DEBIT:0] score_4_x499;
wire signed [DEBIT:0] score_4_x500;
wire signed [DEBIT:0] score_4_x501;
wire signed [DEBIT:0] score_4_x502;
wire signed [DEBIT:0] score_4_x503;
wire signed [DEBIT:0] score_4_x504;
wire signed [DEBIT:0] score_4_x505;
wire signed [DEBIT:0] score_4_x506;
wire signed [DEBIT:0] score_4_x507;
wire signed [DEBIT:0] score_4_x508;
wire signed [DEBIT:0] score_4_x509;
wire signed [DEBIT:0] score_4_x510;
wire signed [DEBIT:0] score_4_x511;
wire signed [DEBIT:0] score_4_x512;
wire signed [DEBIT:0] score_4_x513;
wire signed [DEBIT:0] score_4_x514;
wire signed [DEBIT:0] score_4_x515;
wire signed [DEBIT:0] score_4_x516;
wire signed [DEBIT:0] score_4_x517;
wire signed [DEBIT:0] score_4_x518;
wire signed [DEBIT:0] score_4_x519;
wire signed [DEBIT:0] score_4_x520;
wire signed [DEBIT:0] score_4_x521;
wire signed [DEBIT:0] score_4_x522;
wire signed [DEBIT:0] score_4_x523;
wire signed [DEBIT:0] score_4_x524;
wire signed [DEBIT:0] score_4_x525;
wire signed [DEBIT:0] score_4_x526;
wire signed [DEBIT:0] score_4_x527;
wire signed [DEBIT:0] score_4_x528;
wire signed [DEBIT:0] score_4_x529;
wire signed [DEBIT:0] score_4_x530;
wire signed [DEBIT:0] score_4_x531;
wire signed [DEBIT:0] score_4_x532;
wire signed [DEBIT:0] score_4_x533;
wire signed [DEBIT:0] score_4_x534;
wire signed [DEBIT:0] score_4_x535;
wire signed [DEBIT:0] score_4_x536;
wire signed [DEBIT:0] score_4_x537;
wire signed [DEBIT:0] score_4_x538;
wire signed [DEBIT:0] score_4_x539;
wire signed [DEBIT:0] score_4_x540;
wire signed [DEBIT:0] score_4_x541;
wire signed [DEBIT:0] score_4_x542;
wire signed [DEBIT:0] score_4_x543;
wire signed [DEBIT:0] score_4_x544;
wire signed [DEBIT:0] score_4_x545;
wire signed [DEBIT:0] score_4_x546;
wire signed [DEBIT:0] score_4_x547;
wire signed [DEBIT:0] score_4_x548;
wire signed [DEBIT:0] score_4_x549;
wire signed [DEBIT:0] score_4_x550;
wire signed [DEBIT:0] score_4_x551;
wire signed [DEBIT:0] score_4_x552;
wire signed [DEBIT:0] score_4_x553;
wire signed [DEBIT:0] score_4_x554;
wire signed [DEBIT:0] score_4_x555;
wire signed [DEBIT:0] score_4_x556;
wire signed [DEBIT:0] score_4_x557;
wire signed [DEBIT:0] score_4_x558;
wire signed [DEBIT:0] score_4_x559;
wire signed [DEBIT:0] score_4_x560;
wire signed [DEBIT:0] score_4_x561;
wire signed [DEBIT:0] score_4_x562;
wire signed [DEBIT:0] score_4_x563;
wire signed [DEBIT:0] score_4_x564;
wire signed [DEBIT:0] score_4_x565;
wire signed [DEBIT:0] score_4_x566;
wire signed [DEBIT:0] score_4_x567;
wire signed [DEBIT:0] score_4_x568;
wire signed [DEBIT:0] score_4_x569;
wire signed [DEBIT:0] score_4_x570;
wire signed [DEBIT:0] score_4_x571;
wire signed [DEBIT:0] score_4_x572;
wire signed [DEBIT:0] score_4_x573;
wire signed [DEBIT:0] score_4_x574;
wire signed [DEBIT:0] score_4_x575;
wire signed [DEBIT:0] score_4_x576;
wire signed [DEBIT:0] score_4_x577;
wire signed [DEBIT:0] score_4_x578;
wire signed [DEBIT:0] score_4_x579;
wire signed [DEBIT:0] score_4_x580;
wire signed [DEBIT:0] score_4_x581;
wire signed [DEBIT:0] score_4_x582;
wire signed [DEBIT:0] score_4_x583;
wire signed [DEBIT:0] score_4_x584;
wire signed [DEBIT:0] score_4_x585;
wire signed [DEBIT:0] score_4_x586;
wire signed [DEBIT:0] score_4_x587;
wire signed [DEBIT:0] score_4_x588;
wire signed [DEBIT:0] score_4_x589;
wire signed [DEBIT:0] score_4_x590;
wire signed [DEBIT:0] score_4_x591;
wire signed [DEBIT:0] score_4_x592;
wire signed [DEBIT:0] score_4_x593;
wire signed [DEBIT:0] score_4_x594;
wire signed [DEBIT:0] score_4_x595;
wire signed [DEBIT:0] score_4_x596;
wire signed [DEBIT:0] score_4_x597;
wire signed [DEBIT:0] score_4_x598;
wire signed [DEBIT:0] score_4_x599;
wire signed [DEBIT:0] score_4_x600;
wire signed [DEBIT:0] score_4_x601;
wire signed [DEBIT:0] score_4_x602;
wire signed [DEBIT:0] score_4_x603;
wire signed [DEBIT:0] score_4_x604;
wire signed [DEBIT:0] score_4_x605;
wire signed [DEBIT:0] score_4_x606;
wire signed [DEBIT:0] score_4_x607;
wire signed [DEBIT:0] score_4_x608;
wire signed [DEBIT:0] score_4_x609;
wire signed [DEBIT:0] score_4_x610;
wire signed [DEBIT:0] score_4_x611;
wire signed [DEBIT:0] score_4_x612;
wire signed [DEBIT:0] score_4_x613;
wire signed [DEBIT:0] score_4_x614;
wire signed [DEBIT:0] score_4_x615;
wire signed [DEBIT:0] score_4_x616;
wire signed [DEBIT:0] score_4_x617;
wire signed [DEBIT:0] score_4_x618;
wire signed [DEBIT:0] score_4_x619;
wire signed [DEBIT:0] score_4_x620;
wire signed [DEBIT:0] score_4_x621;
wire signed [DEBIT:0] score_4_x622;
wire signed [DEBIT:0] score_4_x623;
wire signed [DEBIT:0] score_4_x624;
wire signed [DEBIT:0] score_4_x625;
wire signed [DEBIT:0] score_4_x626;
wire signed [DEBIT:0] score_4_x627;
wire signed [DEBIT:0] score_4_x628;
wire signed [DEBIT:0] score_4_x629;
wire signed [DEBIT:0] score_4_x630;
wire signed [DEBIT:0] score_4_x631;
wire signed [DEBIT:0] score_4_x632;
wire signed [DEBIT:0] score_4_x633;
wire signed [DEBIT:0] score_4_x634;
wire signed [DEBIT:0] score_4_x635;
wire signed [DEBIT:0] score_4_x636;
wire signed [DEBIT:0] score_4_x637;
wire signed [DEBIT:0] score_4_x638;
wire signed [DEBIT:0] score_4_x639;
wire signed [DEBIT:0] score_4_x640;
wire signed [DEBIT:0] score_4_x641;
wire signed [DEBIT:0] score_4_x642;
wire signed [DEBIT:0] score_4_x643;
wire signed [DEBIT:0] score_4_x644;
wire signed [DEBIT:0] score_4_x645;
wire signed [DEBIT:0] score_4_x646;
wire signed [DEBIT:0] score_4_x647;
wire signed [DEBIT:0] score_4_x648;
wire signed [DEBIT:0] score_4_x649;
wire signed [DEBIT:0] score_4_x650;
wire signed [DEBIT:0] score_4_x651;
wire signed [DEBIT:0] score_4_x652;
wire signed [DEBIT:0] score_4_x653;
wire signed [DEBIT:0] score_4_x654;
wire signed [DEBIT:0] score_4_x655;
wire signed [DEBIT:0] score_4_x656;
wire signed [DEBIT:0] score_4_x657;
wire signed [DEBIT:0] score_4_x658;
wire signed [DEBIT:0] score_4_x659;
wire signed [DEBIT:0] score_4_x660;
wire signed [DEBIT:0] score_4_x661;
wire signed [DEBIT:0] score_4_x662;
wire signed [DEBIT:0] score_4_x663;
wire signed [DEBIT:0] score_4_x664;
wire signed [DEBIT:0] score_4_x665;
wire signed [DEBIT:0] score_4_x666;
wire signed [DEBIT:0] score_4_x667;
wire signed [DEBIT:0] score_4_x668;
wire signed [DEBIT:0] score_4_x669;
wire signed [DEBIT:0] score_4_x670;
wire signed [DEBIT:0] score_4_x671;
wire signed [DEBIT:0] score_4_x672;
wire signed [DEBIT:0] score_4_x673;
wire signed [DEBIT:0] score_4_x674;
wire signed [DEBIT:0] score_4_x675;
wire signed [DEBIT:0] score_4_x676;
wire signed [DEBIT:0] score_4_x677;
wire signed [DEBIT:0] score_4_x678;
wire signed [DEBIT:0] score_4_x679;
wire signed [DEBIT:0] score_4_x680;
wire signed [DEBIT:0] score_4_x681;
wire signed [DEBIT:0] score_4_x682;
wire signed [DEBIT:0] score_4_x683;
wire signed [DEBIT:0] score_4_x684;
wire signed [DEBIT:0] score_4_x685;
wire signed [DEBIT:0] score_4_x686;
wire signed [DEBIT:0] score_4_x687;
wire signed [DEBIT:0] score_4_x688;
wire signed [DEBIT:0] score_4_x689;
wire signed [DEBIT:0] score_4_x690;
wire signed [DEBIT:0] score_4_x691;
wire signed [DEBIT:0] score_4_x692;
wire signed [DEBIT:0] score_4_x693;
wire signed [DEBIT:0] score_4_x694;
wire signed [DEBIT:0] score_4_x695;
wire signed [DEBIT:0] score_4_x696;
wire signed [DEBIT:0] score_4_x697;
wire signed [DEBIT:0] score_4_x698;
wire signed [DEBIT:0] score_4_x699;
wire signed [DEBIT:0] score_4_x700;
wire signed [DEBIT:0] score_4_x701;
wire signed [DEBIT:0] score_4_x702;
wire signed [DEBIT:0] score_4_x703;
wire signed [DEBIT:0] score_4_x704;
wire signed [DEBIT:0] score_4_x705;
wire signed [DEBIT:0] score_4_x706;
wire signed [DEBIT:0] score_4_x707;
wire signed [DEBIT:0] score_4_x708;
wire signed [DEBIT:0] score_4_x709;
wire signed [DEBIT:0] score_4_x710;
wire signed [DEBIT:0] score_4_x711;
wire signed [DEBIT:0] score_4_x712;
wire signed [DEBIT:0] score_4_x713;
wire signed [DEBIT:0] score_4_x714;
wire signed [DEBIT:0] score_4_x715;
wire signed [DEBIT:0] score_4_x716;
wire signed [DEBIT:0] score_4_x717;
wire signed [DEBIT:0] score_4_x718;
wire signed [DEBIT:0] score_4_x719;
wire signed [DEBIT:0] score_4_x720;
wire signed [DEBIT:0] score_4_x721;
wire signed [DEBIT:0] score_4_x722;
wire signed [DEBIT:0] score_4_x723;
wire signed [DEBIT:0] score_4_x724;
wire signed [DEBIT:0] score_4_x725;
wire signed [DEBIT:0] score_4_x726;
wire signed [DEBIT:0] score_4_x727;
wire signed [DEBIT:0] score_4_x728;
wire signed [DEBIT:0] score_4_x729;
wire signed [DEBIT:0] score_4_x730;
wire signed [DEBIT:0] score_4_x731;
wire signed [DEBIT:0] score_4_x732;
wire signed [DEBIT:0] score_4_x733;
wire signed [DEBIT:0] score_4_x734;
wire signed [DEBIT:0] score_4_x735;
wire signed [DEBIT:0] score_4_x736;
wire signed [DEBIT:0] score_4_x737;
wire signed [DEBIT:0] score_4_x738;
wire signed [DEBIT:0] score_4_x739;
wire signed [DEBIT:0] score_4_x740;
wire signed [DEBIT:0] score_4_x741;
wire signed [DEBIT:0] score_4_x742;
wire signed [DEBIT:0] score_4_x743;
wire signed [DEBIT:0] score_4_x744;
wire signed [DEBIT:0] score_4_x745;
wire signed [DEBIT:0] score_4_x746;
wire signed [DEBIT:0] score_4_x747;
wire signed [DEBIT:0] score_4_x748;
wire signed [DEBIT:0] score_4_x749;
wire signed [DEBIT:0] score_4_x750;
wire signed [DEBIT:0] score_4_x751;
wire signed [DEBIT:0] score_4_x752;
wire signed [DEBIT:0] score_4_x753;
wire signed [DEBIT:0] score_4_x754;
wire signed [DEBIT:0] score_4_x755;
wire signed [DEBIT:0] score_4_x756;
wire signed [DEBIT:0] score_4_x757;
wire signed [DEBIT:0] score_4_x758;
wire signed [DEBIT:0] score_4_x759;
wire signed [DEBIT:0] score_4_x760;
wire signed [DEBIT:0] score_4_x761;
wire signed [DEBIT:0] score_4_x762;
wire signed [DEBIT:0] score_4_x763;
wire signed [DEBIT:0] score_4_x764;
wire signed [DEBIT:0] score_4_x765;
wire signed [DEBIT:0] score_4_x766;
wire signed [DEBIT:0] score_4_x767;
wire signed [DEBIT:0] score_4_x768;
wire signed [DEBIT:0] score_4_x769;
wire signed [DEBIT:0] score_4_x770;
wire signed [DEBIT:0] score_4_x771;
wire signed [DEBIT:0] score_4_x772;
wire signed [DEBIT:0] score_4_x773;
wire signed [DEBIT:0] score_4_x774;
wire signed [DEBIT:0] score_4_x775;
wire signed [DEBIT:0] score_4_x776;
wire signed [DEBIT:0] score_4_x777;
wire signed [DEBIT:0] score_4_x778;
wire signed [DEBIT:0] score_4_x779;
wire signed [DEBIT:0] score_4_x780;
wire signed [DEBIT:0] score_4_x781;
wire signed [DEBIT:0] score_4_x782;
wire signed [DEBIT:0] score_4_x783;
wire signed [DEBIT:0] score_4_x784;
wire signed [DEBIT:0] score_5_x1;
wire signed [DEBIT:0] score_5_x2;
wire signed [DEBIT:0] score_5_x3;
wire signed [DEBIT:0] score_5_x4;
wire signed [DEBIT:0] score_5_x5;
wire signed [DEBIT:0] score_5_x6;
wire signed [DEBIT:0] score_5_x7;
wire signed [DEBIT:0] score_5_x8;
wire signed [DEBIT:0] score_5_x9;
wire signed [DEBIT:0] score_5_x10;
wire signed [DEBIT:0] score_5_x11;
wire signed [DEBIT:0] score_5_x12;
wire signed [DEBIT:0] score_5_x13;
wire signed [DEBIT:0] score_5_x14;
wire signed [DEBIT:0] score_5_x15;
wire signed [DEBIT:0] score_5_x16;
wire signed [DEBIT:0] score_5_x17;
wire signed [DEBIT:0] score_5_x18;
wire signed [DEBIT:0] score_5_x19;
wire signed [DEBIT:0] score_5_x20;
wire signed [DEBIT:0] score_5_x21;
wire signed [DEBIT:0] score_5_x22;
wire signed [DEBIT:0] score_5_x23;
wire signed [DEBIT:0] score_5_x24;
wire signed [DEBIT:0] score_5_x25;
wire signed [DEBIT:0] score_5_x26;
wire signed [DEBIT:0] score_5_x27;
wire signed [DEBIT:0] score_5_x28;
wire signed [DEBIT:0] score_5_x29;
wire signed [DEBIT:0] score_5_x30;
wire signed [DEBIT:0] score_5_x31;
wire signed [DEBIT:0] score_5_x32;
wire signed [DEBIT:0] score_5_x33;
wire signed [DEBIT:0] score_5_x34;
wire signed [DEBIT:0] score_5_x35;
wire signed [DEBIT:0] score_5_x36;
wire signed [DEBIT:0] score_5_x37;
wire signed [DEBIT:0] score_5_x38;
wire signed [DEBIT:0] score_5_x39;
wire signed [DEBIT:0] score_5_x40;
wire signed [DEBIT:0] score_5_x41;
wire signed [DEBIT:0] score_5_x42;
wire signed [DEBIT:0] score_5_x43;
wire signed [DEBIT:0] score_5_x44;
wire signed [DEBIT:0] score_5_x45;
wire signed [DEBIT:0] score_5_x46;
wire signed [DEBIT:0] score_5_x47;
wire signed [DEBIT:0] score_5_x48;
wire signed [DEBIT:0] score_5_x49;
wire signed [DEBIT:0] score_5_x50;
wire signed [DEBIT:0] score_5_x51;
wire signed [DEBIT:0] score_5_x52;
wire signed [DEBIT:0] score_5_x53;
wire signed [DEBIT:0] score_5_x54;
wire signed [DEBIT:0] score_5_x55;
wire signed [DEBIT:0] score_5_x56;
wire signed [DEBIT:0] score_5_x57;
wire signed [DEBIT:0] score_5_x58;
wire signed [DEBIT:0] score_5_x59;
wire signed [DEBIT:0] score_5_x60;
wire signed [DEBIT:0] score_5_x61;
wire signed [DEBIT:0] score_5_x62;
wire signed [DEBIT:0] score_5_x63;
wire signed [DEBIT:0] score_5_x64;
wire signed [DEBIT:0] score_5_x65;
wire signed [DEBIT:0] score_5_x66;
wire signed [DEBIT:0] score_5_x67;
wire signed [DEBIT:0] score_5_x68;
wire signed [DEBIT:0] score_5_x69;
wire signed [DEBIT:0] score_5_x70;
wire signed [DEBIT:0] score_5_x71;
wire signed [DEBIT:0] score_5_x72;
wire signed [DEBIT:0] score_5_x73;
wire signed [DEBIT:0] score_5_x74;
wire signed [DEBIT:0] score_5_x75;
wire signed [DEBIT:0] score_5_x76;
wire signed [DEBIT:0] score_5_x77;
wire signed [DEBIT:0] score_5_x78;
wire signed [DEBIT:0] score_5_x79;
wire signed [DEBIT:0] score_5_x80;
wire signed [DEBIT:0] score_5_x81;
wire signed [DEBIT:0] score_5_x82;
wire signed [DEBIT:0] score_5_x83;
wire signed [DEBIT:0] score_5_x84;
wire signed [DEBIT:0] score_5_x85;
wire signed [DEBIT:0] score_5_x86;
wire signed [DEBIT:0] score_5_x87;
wire signed [DEBIT:0] score_5_x88;
wire signed [DEBIT:0] score_5_x89;
wire signed [DEBIT:0] score_5_x90;
wire signed [DEBIT:0] score_5_x91;
wire signed [DEBIT:0] score_5_x92;
wire signed [DEBIT:0] score_5_x93;
wire signed [DEBIT:0] score_5_x94;
wire signed [DEBIT:0] score_5_x95;
wire signed [DEBIT:0] score_5_x96;
wire signed [DEBIT:0] score_5_x97;
wire signed [DEBIT:0] score_5_x98;
wire signed [DEBIT:0] score_5_x99;
wire signed [DEBIT:0] score_5_x100;
wire signed [DEBIT:0] score_5_x101;
wire signed [DEBIT:0] score_5_x102;
wire signed [DEBIT:0] score_5_x103;
wire signed [DEBIT:0] score_5_x104;
wire signed [DEBIT:0] score_5_x105;
wire signed [DEBIT:0] score_5_x106;
wire signed [DEBIT:0] score_5_x107;
wire signed [DEBIT:0] score_5_x108;
wire signed [DEBIT:0] score_5_x109;
wire signed [DEBIT:0] score_5_x110;
wire signed [DEBIT:0] score_5_x111;
wire signed [DEBIT:0] score_5_x112;
wire signed [DEBIT:0] score_5_x113;
wire signed [DEBIT:0] score_5_x114;
wire signed [DEBIT:0] score_5_x115;
wire signed [DEBIT:0] score_5_x116;
wire signed [DEBIT:0] score_5_x117;
wire signed [DEBIT:0] score_5_x118;
wire signed [DEBIT:0] score_5_x119;
wire signed [DEBIT:0] score_5_x120;
wire signed [DEBIT:0] score_5_x121;
wire signed [DEBIT:0] score_5_x122;
wire signed [DEBIT:0] score_5_x123;
wire signed [DEBIT:0] score_5_x124;
wire signed [DEBIT:0] score_5_x125;
wire signed [DEBIT:0] score_5_x126;
wire signed [DEBIT:0] score_5_x127;
wire signed [DEBIT:0] score_5_x128;
wire signed [DEBIT:0] score_5_x129;
wire signed [DEBIT:0] score_5_x130;
wire signed [DEBIT:0] score_5_x131;
wire signed [DEBIT:0] score_5_x132;
wire signed [DEBIT:0] score_5_x133;
wire signed [DEBIT:0] score_5_x134;
wire signed [DEBIT:0] score_5_x135;
wire signed [DEBIT:0] score_5_x136;
wire signed [DEBIT:0] score_5_x137;
wire signed [DEBIT:0] score_5_x138;
wire signed [DEBIT:0] score_5_x139;
wire signed [DEBIT:0] score_5_x140;
wire signed [DEBIT:0] score_5_x141;
wire signed [DEBIT:0] score_5_x142;
wire signed [DEBIT:0] score_5_x143;
wire signed [DEBIT:0] score_5_x144;
wire signed [DEBIT:0] score_5_x145;
wire signed [DEBIT:0] score_5_x146;
wire signed [DEBIT:0] score_5_x147;
wire signed [DEBIT:0] score_5_x148;
wire signed [DEBIT:0] score_5_x149;
wire signed [DEBIT:0] score_5_x150;
wire signed [DEBIT:0] score_5_x151;
wire signed [DEBIT:0] score_5_x152;
wire signed [DEBIT:0] score_5_x153;
wire signed [DEBIT:0] score_5_x154;
wire signed [DEBIT:0] score_5_x155;
wire signed [DEBIT:0] score_5_x156;
wire signed [DEBIT:0] score_5_x157;
wire signed [DEBIT:0] score_5_x158;
wire signed [DEBIT:0] score_5_x159;
wire signed [DEBIT:0] score_5_x160;
wire signed [DEBIT:0] score_5_x161;
wire signed [DEBIT:0] score_5_x162;
wire signed [DEBIT:0] score_5_x163;
wire signed [DEBIT:0] score_5_x164;
wire signed [DEBIT:0] score_5_x165;
wire signed [DEBIT:0] score_5_x166;
wire signed [DEBIT:0] score_5_x167;
wire signed [DEBIT:0] score_5_x168;
wire signed [DEBIT:0] score_5_x169;
wire signed [DEBIT:0] score_5_x170;
wire signed [DEBIT:0] score_5_x171;
wire signed [DEBIT:0] score_5_x172;
wire signed [DEBIT:0] score_5_x173;
wire signed [DEBIT:0] score_5_x174;
wire signed [DEBIT:0] score_5_x175;
wire signed [DEBIT:0] score_5_x176;
wire signed [DEBIT:0] score_5_x177;
wire signed [DEBIT:0] score_5_x178;
wire signed [DEBIT:0] score_5_x179;
wire signed [DEBIT:0] score_5_x180;
wire signed [DEBIT:0] score_5_x181;
wire signed [DEBIT:0] score_5_x182;
wire signed [DEBIT:0] score_5_x183;
wire signed [DEBIT:0] score_5_x184;
wire signed [DEBIT:0] score_5_x185;
wire signed [DEBIT:0] score_5_x186;
wire signed [DEBIT:0] score_5_x187;
wire signed [DEBIT:0] score_5_x188;
wire signed [DEBIT:0] score_5_x189;
wire signed [DEBIT:0] score_5_x190;
wire signed [DEBIT:0] score_5_x191;
wire signed [DEBIT:0] score_5_x192;
wire signed [DEBIT:0] score_5_x193;
wire signed [DEBIT:0] score_5_x194;
wire signed [DEBIT:0] score_5_x195;
wire signed [DEBIT:0] score_5_x196;
wire signed [DEBIT:0] score_5_x197;
wire signed [DEBIT:0] score_5_x198;
wire signed [DEBIT:0] score_5_x199;
wire signed [DEBIT:0] score_5_x200;
wire signed [DEBIT:0] score_5_x201;
wire signed [DEBIT:0] score_5_x202;
wire signed [DEBIT:0] score_5_x203;
wire signed [DEBIT:0] score_5_x204;
wire signed [DEBIT:0] score_5_x205;
wire signed [DEBIT:0] score_5_x206;
wire signed [DEBIT:0] score_5_x207;
wire signed [DEBIT:0] score_5_x208;
wire signed [DEBIT:0] score_5_x209;
wire signed [DEBIT:0] score_5_x210;
wire signed [DEBIT:0] score_5_x211;
wire signed [DEBIT:0] score_5_x212;
wire signed [DEBIT:0] score_5_x213;
wire signed [DEBIT:0] score_5_x214;
wire signed [DEBIT:0] score_5_x215;
wire signed [DEBIT:0] score_5_x216;
wire signed [DEBIT:0] score_5_x217;
wire signed [DEBIT:0] score_5_x218;
wire signed [DEBIT:0] score_5_x219;
wire signed [DEBIT:0] score_5_x220;
wire signed [DEBIT:0] score_5_x221;
wire signed [DEBIT:0] score_5_x222;
wire signed [DEBIT:0] score_5_x223;
wire signed [DEBIT:0] score_5_x224;
wire signed [DEBIT:0] score_5_x225;
wire signed [DEBIT:0] score_5_x226;
wire signed [DEBIT:0] score_5_x227;
wire signed [DEBIT:0] score_5_x228;
wire signed [DEBIT:0] score_5_x229;
wire signed [DEBIT:0] score_5_x230;
wire signed [DEBIT:0] score_5_x231;
wire signed [DEBIT:0] score_5_x232;
wire signed [DEBIT:0] score_5_x233;
wire signed [DEBIT:0] score_5_x234;
wire signed [DEBIT:0] score_5_x235;
wire signed [DEBIT:0] score_5_x236;
wire signed [DEBIT:0] score_5_x237;
wire signed [DEBIT:0] score_5_x238;
wire signed [DEBIT:0] score_5_x239;
wire signed [DEBIT:0] score_5_x240;
wire signed [DEBIT:0] score_5_x241;
wire signed [DEBIT:0] score_5_x242;
wire signed [DEBIT:0] score_5_x243;
wire signed [DEBIT:0] score_5_x244;
wire signed [DEBIT:0] score_5_x245;
wire signed [DEBIT:0] score_5_x246;
wire signed [DEBIT:0] score_5_x247;
wire signed [DEBIT:0] score_5_x248;
wire signed [DEBIT:0] score_5_x249;
wire signed [DEBIT:0] score_5_x250;
wire signed [DEBIT:0] score_5_x251;
wire signed [DEBIT:0] score_5_x252;
wire signed [DEBIT:0] score_5_x253;
wire signed [DEBIT:0] score_5_x254;
wire signed [DEBIT:0] score_5_x255;
wire signed [DEBIT:0] score_5_x256;
wire signed [DEBIT:0] score_5_x257;
wire signed [DEBIT:0] score_5_x258;
wire signed [DEBIT:0] score_5_x259;
wire signed [DEBIT:0] score_5_x260;
wire signed [DEBIT:0] score_5_x261;
wire signed [DEBIT:0] score_5_x262;
wire signed [DEBIT:0] score_5_x263;
wire signed [DEBIT:0] score_5_x264;
wire signed [DEBIT:0] score_5_x265;
wire signed [DEBIT:0] score_5_x266;
wire signed [DEBIT:0] score_5_x267;
wire signed [DEBIT:0] score_5_x268;
wire signed [DEBIT:0] score_5_x269;
wire signed [DEBIT:0] score_5_x270;
wire signed [DEBIT:0] score_5_x271;
wire signed [DEBIT:0] score_5_x272;
wire signed [DEBIT:0] score_5_x273;
wire signed [DEBIT:0] score_5_x274;
wire signed [DEBIT:0] score_5_x275;
wire signed [DEBIT:0] score_5_x276;
wire signed [DEBIT:0] score_5_x277;
wire signed [DEBIT:0] score_5_x278;
wire signed [DEBIT:0] score_5_x279;
wire signed [DEBIT:0] score_5_x280;
wire signed [DEBIT:0] score_5_x281;
wire signed [DEBIT:0] score_5_x282;
wire signed [DEBIT:0] score_5_x283;
wire signed [DEBIT:0] score_5_x284;
wire signed [DEBIT:0] score_5_x285;
wire signed [DEBIT:0] score_5_x286;
wire signed [DEBIT:0] score_5_x287;
wire signed [DEBIT:0] score_5_x288;
wire signed [DEBIT:0] score_5_x289;
wire signed [DEBIT:0] score_5_x290;
wire signed [DEBIT:0] score_5_x291;
wire signed [DEBIT:0] score_5_x292;
wire signed [DEBIT:0] score_5_x293;
wire signed [DEBIT:0] score_5_x294;
wire signed [DEBIT:0] score_5_x295;
wire signed [DEBIT:0] score_5_x296;
wire signed [DEBIT:0] score_5_x297;
wire signed [DEBIT:0] score_5_x298;
wire signed [DEBIT:0] score_5_x299;
wire signed [DEBIT:0] score_5_x300;
wire signed [DEBIT:0] score_5_x301;
wire signed [DEBIT:0] score_5_x302;
wire signed [DEBIT:0] score_5_x303;
wire signed [DEBIT:0] score_5_x304;
wire signed [DEBIT:0] score_5_x305;
wire signed [DEBIT:0] score_5_x306;
wire signed [DEBIT:0] score_5_x307;
wire signed [DEBIT:0] score_5_x308;
wire signed [DEBIT:0] score_5_x309;
wire signed [DEBIT:0] score_5_x310;
wire signed [DEBIT:0] score_5_x311;
wire signed [DEBIT:0] score_5_x312;
wire signed [DEBIT:0] score_5_x313;
wire signed [DEBIT:0] score_5_x314;
wire signed [DEBIT:0] score_5_x315;
wire signed [DEBIT:0] score_5_x316;
wire signed [DEBIT:0] score_5_x317;
wire signed [DEBIT:0] score_5_x318;
wire signed [DEBIT:0] score_5_x319;
wire signed [DEBIT:0] score_5_x320;
wire signed [DEBIT:0] score_5_x321;
wire signed [DEBIT:0] score_5_x322;
wire signed [DEBIT:0] score_5_x323;
wire signed [DEBIT:0] score_5_x324;
wire signed [DEBIT:0] score_5_x325;
wire signed [DEBIT:0] score_5_x326;
wire signed [DEBIT:0] score_5_x327;
wire signed [DEBIT:0] score_5_x328;
wire signed [DEBIT:0] score_5_x329;
wire signed [DEBIT:0] score_5_x330;
wire signed [DEBIT:0] score_5_x331;
wire signed [DEBIT:0] score_5_x332;
wire signed [DEBIT:0] score_5_x333;
wire signed [DEBIT:0] score_5_x334;
wire signed [DEBIT:0] score_5_x335;
wire signed [DEBIT:0] score_5_x336;
wire signed [DEBIT:0] score_5_x337;
wire signed [DEBIT:0] score_5_x338;
wire signed [DEBIT:0] score_5_x339;
wire signed [DEBIT:0] score_5_x340;
wire signed [DEBIT:0] score_5_x341;
wire signed [DEBIT:0] score_5_x342;
wire signed [DEBIT:0] score_5_x343;
wire signed [DEBIT:0] score_5_x344;
wire signed [DEBIT:0] score_5_x345;
wire signed [DEBIT:0] score_5_x346;
wire signed [DEBIT:0] score_5_x347;
wire signed [DEBIT:0] score_5_x348;
wire signed [DEBIT:0] score_5_x349;
wire signed [DEBIT:0] score_5_x350;
wire signed [DEBIT:0] score_5_x351;
wire signed [DEBIT:0] score_5_x352;
wire signed [DEBIT:0] score_5_x353;
wire signed [DEBIT:0] score_5_x354;
wire signed [DEBIT:0] score_5_x355;
wire signed [DEBIT:0] score_5_x356;
wire signed [DEBIT:0] score_5_x357;
wire signed [DEBIT:0] score_5_x358;
wire signed [DEBIT:0] score_5_x359;
wire signed [DEBIT:0] score_5_x360;
wire signed [DEBIT:0] score_5_x361;
wire signed [DEBIT:0] score_5_x362;
wire signed [DEBIT:0] score_5_x363;
wire signed [DEBIT:0] score_5_x364;
wire signed [DEBIT:0] score_5_x365;
wire signed [DEBIT:0] score_5_x366;
wire signed [DEBIT:0] score_5_x367;
wire signed [DEBIT:0] score_5_x368;
wire signed [DEBIT:0] score_5_x369;
wire signed [DEBIT:0] score_5_x370;
wire signed [DEBIT:0] score_5_x371;
wire signed [DEBIT:0] score_5_x372;
wire signed [DEBIT:0] score_5_x373;
wire signed [DEBIT:0] score_5_x374;
wire signed [DEBIT:0] score_5_x375;
wire signed [DEBIT:0] score_5_x376;
wire signed [DEBIT:0] score_5_x377;
wire signed [DEBIT:0] score_5_x378;
wire signed [DEBIT:0] score_5_x379;
wire signed [DEBIT:0] score_5_x380;
wire signed [DEBIT:0] score_5_x381;
wire signed [DEBIT:0] score_5_x382;
wire signed [DEBIT:0] score_5_x383;
wire signed [DEBIT:0] score_5_x384;
wire signed [DEBIT:0] score_5_x385;
wire signed [DEBIT:0] score_5_x386;
wire signed [DEBIT:0] score_5_x387;
wire signed [DEBIT:0] score_5_x388;
wire signed [DEBIT:0] score_5_x389;
wire signed [DEBIT:0] score_5_x390;
wire signed [DEBIT:0] score_5_x391;
wire signed [DEBIT:0] score_5_x392;
wire signed [DEBIT:0] score_5_x393;
wire signed [DEBIT:0] score_5_x394;
wire signed [DEBIT:0] score_5_x395;
wire signed [DEBIT:0] score_5_x396;
wire signed [DEBIT:0] score_5_x397;
wire signed [DEBIT:0] score_5_x398;
wire signed [DEBIT:0] score_5_x399;
wire signed [DEBIT:0] score_5_x400;
wire signed [DEBIT:0] score_5_x401;
wire signed [DEBIT:0] score_5_x402;
wire signed [DEBIT:0] score_5_x403;
wire signed [DEBIT:0] score_5_x404;
wire signed [DEBIT:0] score_5_x405;
wire signed [DEBIT:0] score_5_x406;
wire signed [DEBIT:0] score_5_x407;
wire signed [DEBIT:0] score_5_x408;
wire signed [DEBIT:0] score_5_x409;
wire signed [DEBIT:0] score_5_x410;
wire signed [DEBIT:0] score_5_x411;
wire signed [DEBIT:0] score_5_x412;
wire signed [DEBIT:0] score_5_x413;
wire signed [DEBIT:0] score_5_x414;
wire signed [DEBIT:0] score_5_x415;
wire signed [DEBIT:0] score_5_x416;
wire signed [DEBIT:0] score_5_x417;
wire signed [DEBIT:0] score_5_x418;
wire signed [DEBIT:0] score_5_x419;
wire signed [DEBIT:0] score_5_x420;
wire signed [DEBIT:0] score_5_x421;
wire signed [DEBIT:0] score_5_x422;
wire signed [DEBIT:0] score_5_x423;
wire signed [DEBIT:0] score_5_x424;
wire signed [DEBIT:0] score_5_x425;
wire signed [DEBIT:0] score_5_x426;
wire signed [DEBIT:0] score_5_x427;
wire signed [DEBIT:0] score_5_x428;
wire signed [DEBIT:0] score_5_x429;
wire signed [DEBIT:0] score_5_x430;
wire signed [DEBIT:0] score_5_x431;
wire signed [DEBIT:0] score_5_x432;
wire signed [DEBIT:0] score_5_x433;
wire signed [DEBIT:0] score_5_x434;
wire signed [DEBIT:0] score_5_x435;
wire signed [DEBIT:0] score_5_x436;
wire signed [DEBIT:0] score_5_x437;
wire signed [DEBIT:0] score_5_x438;
wire signed [DEBIT:0] score_5_x439;
wire signed [DEBIT:0] score_5_x440;
wire signed [DEBIT:0] score_5_x441;
wire signed [DEBIT:0] score_5_x442;
wire signed [DEBIT:0] score_5_x443;
wire signed [DEBIT:0] score_5_x444;
wire signed [DEBIT:0] score_5_x445;
wire signed [DEBIT:0] score_5_x446;
wire signed [DEBIT:0] score_5_x447;
wire signed [DEBIT:0] score_5_x448;
wire signed [DEBIT:0] score_5_x449;
wire signed [DEBIT:0] score_5_x450;
wire signed [DEBIT:0] score_5_x451;
wire signed [DEBIT:0] score_5_x452;
wire signed [DEBIT:0] score_5_x453;
wire signed [DEBIT:0] score_5_x454;
wire signed [DEBIT:0] score_5_x455;
wire signed [DEBIT:0] score_5_x456;
wire signed [DEBIT:0] score_5_x457;
wire signed [DEBIT:0] score_5_x458;
wire signed [DEBIT:0] score_5_x459;
wire signed [DEBIT:0] score_5_x460;
wire signed [DEBIT:0] score_5_x461;
wire signed [DEBIT:0] score_5_x462;
wire signed [DEBIT:0] score_5_x463;
wire signed [DEBIT:0] score_5_x464;
wire signed [DEBIT:0] score_5_x465;
wire signed [DEBIT:0] score_5_x466;
wire signed [DEBIT:0] score_5_x467;
wire signed [DEBIT:0] score_5_x468;
wire signed [DEBIT:0] score_5_x469;
wire signed [DEBIT:0] score_5_x470;
wire signed [DEBIT:0] score_5_x471;
wire signed [DEBIT:0] score_5_x472;
wire signed [DEBIT:0] score_5_x473;
wire signed [DEBIT:0] score_5_x474;
wire signed [DEBIT:0] score_5_x475;
wire signed [DEBIT:0] score_5_x476;
wire signed [DEBIT:0] score_5_x477;
wire signed [DEBIT:0] score_5_x478;
wire signed [DEBIT:0] score_5_x479;
wire signed [DEBIT:0] score_5_x480;
wire signed [DEBIT:0] score_5_x481;
wire signed [DEBIT:0] score_5_x482;
wire signed [DEBIT:0] score_5_x483;
wire signed [DEBIT:0] score_5_x484;
wire signed [DEBIT:0] score_5_x485;
wire signed [DEBIT:0] score_5_x486;
wire signed [DEBIT:0] score_5_x487;
wire signed [DEBIT:0] score_5_x488;
wire signed [DEBIT:0] score_5_x489;
wire signed [DEBIT:0] score_5_x490;
wire signed [DEBIT:0] score_5_x491;
wire signed [DEBIT:0] score_5_x492;
wire signed [DEBIT:0] score_5_x493;
wire signed [DEBIT:0] score_5_x494;
wire signed [DEBIT:0] score_5_x495;
wire signed [DEBIT:0] score_5_x496;
wire signed [DEBIT:0] score_5_x497;
wire signed [DEBIT:0] score_5_x498;
wire signed [DEBIT:0] score_5_x499;
wire signed [DEBIT:0] score_5_x500;
wire signed [DEBIT:0] score_5_x501;
wire signed [DEBIT:0] score_5_x502;
wire signed [DEBIT:0] score_5_x503;
wire signed [DEBIT:0] score_5_x504;
wire signed [DEBIT:0] score_5_x505;
wire signed [DEBIT:0] score_5_x506;
wire signed [DEBIT:0] score_5_x507;
wire signed [DEBIT:0] score_5_x508;
wire signed [DEBIT:0] score_5_x509;
wire signed [DEBIT:0] score_5_x510;
wire signed [DEBIT:0] score_5_x511;
wire signed [DEBIT:0] score_5_x512;
wire signed [DEBIT:0] score_5_x513;
wire signed [DEBIT:0] score_5_x514;
wire signed [DEBIT:0] score_5_x515;
wire signed [DEBIT:0] score_5_x516;
wire signed [DEBIT:0] score_5_x517;
wire signed [DEBIT:0] score_5_x518;
wire signed [DEBIT:0] score_5_x519;
wire signed [DEBIT:0] score_5_x520;
wire signed [DEBIT:0] score_5_x521;
wire signed [DEBIT:0] score_5_x522;
wire signed [DEBIT:0] score_5_x523;
wire signed [DEBIT:0] score_5_x524;
wire signed [DEBIT:0] score_5_x525;
wire signed [DEBIT:0] score_5_x526;
wire signed [DEBIT:0] score_5_x527;
wire signed [DEBIT:0] score_5_x528;
wire signed [DEBIT:0] score_5_x529;
wire signed [DEBIT:0] score_5_x530;
wire signed [DEBIT:0] score_5_x531;
wire signed [DEBIT:0] score_5_x532;
wire signed [DEBIT:0] score_5_x533;
wire signed [DEBIT:0] score_5_x534;
wire signed [DEBIT:0] score_5_x535;
wire signed [DEBIT:0] score_5_x536;
wire signed [DEBIT:0] score_5_x537;
wire signed [DEBIT:0] score_5_x538;
wire signed [DEBIT:0] score_5_x539;
wire signed [DEBIT:0] score_5_x540;
wire signed [DEBIT:0] score_5_x541;
wire signed [DEBIT:0] score_5_x542;
wire signed [DEBIT:0] score_5_x543;
wire signed [DEBIT:0] score_5_x544;
wire signed [DEBIT:0] score_5_x545;
wire signed [DEBIT:0] score_5_x546;
wire signed [DEBIT:0] score_5_x547;
wire signed [DEBIT:0] score_5_x548;
wire signed [DEBIT:0] score_5_x549;
wire signed [DEBIT:0] score_5_x550;
wire signed [DEBIT:0] score_5_x551;
wire signed [DEBIT:0] score_5_x552;
wire signed [DEBIT:0] score_5_x553;
wire signed [DEBIT:0] score_5_x554;
wire signed [DEBIT:0] score_5_x555;
wire signed [DEBIT:0] score_5_x556;
wire signed [DEBIT:0] score_5_x557;
wire signed [DEBIT:0] score_5_x558;
wire signed [DEBIT:0] score_5_x559;
wire signed [DEBIT:0] score_5_x560;
wire signed [DEBIT:0] score_5_x561;
wire signed [DEBIT:0] score_5_x562;
wire signed [DEBIT:0] score_5_x563;
wire signed [DEBIT:0] score_5_x564;
wire signed [DEBIT:0] score_5_x565;
wire signed [DEBIT:0] score_5_x566;
wire signed [DEBIT:0] score_5_x567;
wire signed [DEBIT:0] score_5_x568;
wire signed [DEBIT:0] score_5_x569;
wire signed [DEBIT:0] score_5_x570;
wire signed [DEBIT:0] score_5_x571;
wire signed [DEBIT:0] score_5_x572;
wire signed [DEBIT:0] score_5_x573;
wire signed [DEBIT:0] score_5_x574;
wire signed [DEBIT:0] score_5_x575;
wire signed [DEBIT:0] score_5_x576;
wire signed [DEBIT:0] score_5_x577;
wire signed [DEBIT:0] score_5_x578;
wire signed [DEBIT:0] score_5_x579;
wire signed [DEBIT:0] score_5_x580;
wire signed [DEBIT:0] score_5_x581;
wire signed [DEBIT:0] score_5_x582;
wire signed [DEBIT:0] score_5_x583;
wire signed [DEBIT:0] score_5_x584;
wire signed [DEBIT:0] score_5_x585;
wire signed [DEBIT:0] score_5_x586;
wire signed [DEBIT:0] score_5_x587;
wire signed [DEBIT:0] score_5_x588;
wire signed [DEBIT:0] score_5_x589;
wire signed [DEBIT:0] score_5_x590;
wire signed [DEBIT:0] score_5_x591;
wire signed [DEBIT:0] score_5_x592;
wire signed [DEBIT:0] score_5_x593;
wire signed [DEBIT:0] score_5_x594;
wire signed [DEBIT:0] score_5_x595;
wire signed [DEBIT:0] score_5_x596;
wire signed [DEBIT:0] score_5_x597;
wire signed [DEBIT:0] score_5_x598;
wire signed [DEBIT:0] score_5_x599;
wire signed [DEBIT:0] score_5_x600;
wire signed [DEBIT:0] score_5_x601;
wire signed [DEBIT:0] score_5_x602;
wire signed [DEBIT:0] score_5_x603;
wire signed [DEBIT:0] score_5_x604;
wire signed [DEBIT:0] score_5_x605;
wire signed [DEBIT:0] score_5_x606;
wire signed [DEBIT:0] score_5_x607;
wire signed [DEBIT:0] score_5_x608;
wire signed [DEBIT:0] score_5_x609;
wire signed [DEBIT:0] score_5_x610;
wire signed [DEBIT:0] score_5_x611;
wire signed [DEBIT:0] score_5_x612;
wire signed [DEBIT:0] score_5_x613;
wire signed [DEBIT:0] score_5_x614;
wire signed [DEBIT:0] score_5_x615;
wire signed [DEBIT:0] score_5_x616;
wire signed [DEBIT:0] score_5_x617;
wire signed [DEBIT:0] score_5_x618;
wire signed [DEBIT:0] score_5_x619;
wire signed [DEBIT:0] score_5_x620;
wire signed [DEBIT:0] score_5_x621;
wire signed [DEBIT:0] score_5_x622;
wire signed [DEBIT:0] score_5_x623;
wire signed [DEBIT:0] score_5_x624;
wire signed [DEBIT:0] score_5_x625;
wire signed [DEBIT:0] score_5_x626;
wire signed [DEBIT:0] score_5_x627;
wire signed [DEBIT:0] score_5_x628;
wire signed [DEBIT:0] score_5_x629;
wire signed [DEBIT:0] score_5_x630;
wire signed [DEBIT:0] score_5_x631;
wire signed [DEBIT:0] score_5_x632;
wire signed [DEBIT:0] score_5_x633;
wire signed [DEBIT:0] score_5_x634;
wire signed [DEBIT:0] score_5_x635;
wire signed [DEBIT:0] score_5_x636;
wire signed [DEBIT:0] score_5_x637;
wire signed [DEBIT:0] score_5_x638;
wire signed [DEBIT:0] score_5_x639;
wire signed [DEBIT:0] score_5_x640;
wire signed [DEBIT:0] score_5_x641;
wire signed [DEBIT:0] score_5_x642;
wire signed [DEBIT:0] score_5_x643;
wire signed [DEBIT:0] score_5_x644;
wire signed [DEBIT:0] score_5_x645;
wire signed [DEBIT:0] score_5_x646;
wire signed [DEBIT:0] score_5_x647;
wire signed [DEBIT:0] score_5_x648;
wire signed [DEBIT:0] score_5_x649;
wire signed [DEBIT:0] score_5_x650;
wire signed [DEBIT:0] score_5_x651;
wire signed [DEBIT:0] score_5_x652;
wire signed [DEBIT:0] score_5_x653;
wire signed [DEBIT:0] score_5_x654;
wire signed [DEBIT:0] score_5_x655;
wire signed [DEBIT:0] score_5_x656;
wire signed [DEBIT:0] score_5_x657;
wire signed [DEBIT:0] score_5_x658;
wire signed [DEBIT:0] score_5_x659;
wire signed [DEBIT:0] score_5_x660;
wire signed [DEBIT:0] score_5_x661;
wire signed [DEBIT:0] score_5_x662;
wire signed [DEBIT:0] score_5_x663;
wire signed [DEBIT:0] score_5_x664;
wire signed [DEBIT:0] score_5_x665;
wire signed [DEBIT:0] score_5_x666;
wire signed [DEBIT:0] score_5_x667;
wire signed [DEBIT:0] score_5_x668;
wire signed [DEBIT:0] score_5_x669;
wire signed [DEBIT:0] score_5_x670;
wire signed [DEBIT:0] score_5_x671;
wire signed [DEBIT:0] score_5_x672;
wire signed [DEBIT:0] score_5_x673;
wire signed [DEBIT:0] score_5_x674;
wire signed [DEBIT:0] score_5_x675;
wire signed [DEBIT:0] score_5_x676;
wire signed [DEBIT:0] score_5_x677;
wire signed [DEBIT:0] score_5_x678;
wire signed [DEBIT:0] score_5_x679;
wire signed [DEBIT:0] score_5_x680;
wire signed [DEBIT:0] score_5_x681;
wire signed [DEBIT:0] score_5_x682;
wire signed [DEBIT:0] score_5_x683;
wire signed [DEBIT:0] score_5_x684;
wire signed [DEBIT:0] score_5_x685;
wire signed [DEBIT:0] score_5_x686;
wire signed [DEBIT:0] score_5_x687;
wire signed [DEBIT:0] score_5_x688;
wire signed [DEBIT:0] score_5_x689;
wire signed [DEBIT:0] score_5_x690;
wire signed [DEBIT:0] score_5_x691;
wire signed [DEBIT:0] score_5_x692;
wire signed [DEBIT:0] score_5_x693;
wire signed [DEBIT:0] score_5_x694;
wire signed [DEBIT:0] score_5_x695;
wire signed [DEBIT:0] score_5_x696;
wire signed [DEBIT:0] score_5_x697;
wire signed [DEBIT:0] score_5_x698;
wire signed [DEBIT:0] score_5_x699;
wire signed [DEBIT:0] score_5_x700;
wire signed [DEBIT:0] score_5_x701;
wire signed [DEBIT:0] score_5_x702;
wire signed [DEBIT:0] score_5_x703;
wire signed [DEBIT:0] score_5_x704;
wire signed [DEBIT:0] score_5_x705;
wire signed [DEBIT:0] score_5_x706;
wire signed [DEBIT:0] score_5_x707;
wire signed [DEBIT:0] score_5_x708;
wire signed [DEBIT:0] score_5_x709;
wire signed [DEBIT:0] score_5_x710;
wire signed [DEBIT:0] score_5_x711;
wire signed [DEBIT:0] score_5_x712;
wire signed [DEBIT:0] score_5_x713;
wire signed [DEBIT:0] score_5_x714;
wire signed [DEBIT:0] score_5_x715;
wire signed [DEBIT:0] score_5_x716;
wire signed [DEBIT:0] score_5_x717;
wire signed [DEBIT:0] score_5_x718;
wire signed [DEBIT:0] score_5_x719;
wire signed [DEBIT:0] score_5_x720;
wire signed [DEBIT:0] score_5_x721;
wire signed [DEBIT:0] score_5_x722;
wire signed [DEBIT:0] score_5_x723;
wire signed [DEBIT:0] score_5_x724;
wire signed [DEBIT:0] score_5_x725;
wire signed [DEBIT:0] score_5_x726;
wire signed [DEBIT:0] score_5_x727;
wire signed [DEBIT:0] score_5_x728;
wire signed [DEBIT:0] score_5_x729;
wire signed [DEBIT:0] score_5_x730;
wire signed [DEBIT:0] score_5_x731;
wire signed [DEBIT:0] score_5_x732;
wire signed [DEBIT:0] score_5_x733;
wire signed [DEBIT:0] score_5_x734;
wire signed [DEBIT:0] score_5_x735;
wire signed [DEBIT:0] score_5_x736;
wire signed [DEBIT:0] score_5_x737;
wire signed [DEBIT:0] score_5_x738;
wire signed [DEBIT:0] score_5_x739;
wire signed [DEBIT:0] score_5_x740;
wire signed [DEBIT:0] score_5_x741;
wire signed [DEBIT:0] score_5_x742;
wire signed [DEBIT:0] score_5_x743;
wire signed [DEBIT:0] score_5_x744;
wire signed [DEBIT:0] score_5_x745;
wire signed [DEBIT:0] score_5_x746;
wire signed [DEBIT:0] score_5_x747;
wire signed [DEBIT:0] score_5_x748;
wire signed [DEBIT:0] score_5_x749;
wire signed [DEBIT:0] score_5_x750;
wire signed [DEBIT:0] score_5_x751;
wire signed [DEBIT:0] score_5_x752;
wire signed [DEBIT:0] score_5_x753;
wire signed [DEBIT:0] score_5_x754;
wire signed [DEBIT:0] score_5_x755;
wire signed [DEBIT:0] score_5_x756;
wire signed [DEBIT:0] score_5_x757;
wire signed [DEBIT:0] score_5_x758;
wire signed [DEBIT:0] score_5_x759;
wire signed [DEBIT:0] score_5_x760;
wire signed [DEBIT:0] score_5_x761;
wire signed [DEBIT:0] score_5_x762;
wire signed [DEBIT:0] score_5_x763;
wire signed [DEBIT:0] score_5_x764;
wire signed [DEBIT:0] score_5_x765;
wire signed [DEBIT:0] score_5_x766;
wire signed [DEBIT:0] score_5_x767;
wire signed [DEBIT:0] score_5_x768;
wire signed [DEBIT:0] score_5_x769;
wire signed [DEBIT:0] score_5_x770;
wire signed [DEBIT:0] score_5_x771;
wire signed [DEBIT:0] score_5_x772;
wire signed [DEBIT:0] score_5_x773;
wire signed [DEBIT:0] score_5_x774;
wire signed [DEBIT:0] score_5_x775;
wire signed [DEBIT:0] score_5_x776;
wire signed [DEBIT:0] score_5_x777;
wire signed [DEBIT:0] score_5_x778;
wire signed [DEBIT:0] score_5_x779;
wire signed [DEBIT:0] score_5_x780;
wire signed [DEBIT:0] score_5_x781;
wire signed [DEBIT:0] score_5_x782;
wire signed [DEBIT:0] score_5_x783;
wire signed [DEBIT:0] score_5_x784;
wire signed [DEBIT:0] score_6_x1;
wire signed [DEBIT:0] score_6_x2;
wire signed [DEBIT:0] score_6_x3;
wire signed [DEBIT:0] score_6_x4;
wire signed [DEBIT:0] score_6_x5;
wire signed [DEBIT:0] score_6_x6;
wire signed [DEBIT:0] score_6_x7;
wire signed [DEBIT:0] score_6_x8;
wire signed [DEBIT:0] score_6_x9;
wire signed [DEBIT:0] score_6_x10;
wire signed [DEBIT:0] score_6_x11;
wire signed [DEBIT:0] score_6_x12;
wire signed [DEBIT:0] score_6_x13;
wire signed [DEBIT:0] score_6_x14;
wire signed [DEBIT:0] score_6_x15;
wire signed [DEBIT:0] score_6_x16;
wire signed [DEBIT:0] score_6_x17;
wire signed [DEBIT:0] score_6_x18;
wire signed [DEBIT:0] score_6_x19;
wire signed [DEBIT:0] score_6_x20;
wire signed [DEBIT:0] score_6_x21;
wire signed [DEBIT:0] score_6_x22;
wire signed [DEBIT:0] score_6_x23;
wire signed [DEBIT:0] score_6_x24;
wire signed [DEBIT:0] score_6_x25;
wire signed [DEBIT:0] score_6_x26;
wire signed [DEBIT:0] score_6_x27;
wire signed [DEBIT:0] score_6_x28;
wire signed [DEBIT:0] score_6_x29;
wire signed [DEBIT:0] score_6_x30;
wire signed [DEBIT:0] score_6_x31;
wire signed [DEBIT:0] score_6_x32;
wire signed [DEBIT:0] score_6_x33;
wire signed [DEBIT:0] score_6_x34;
wire signed [DEBIT:0] score_6_x35;
wire signed [DEBIT:0] score_6_x36;
wire signed [DEBIT:0] score_6_x37;
wire signed [DEBIT:0] score_6_x38;
wire signed [DEBIT:0] score_6_x39;
wire signed [DEBIT:0] score_6_x40;
wire signed [DEBIT:0] score_6_x41;
wire signed [DEBIT:0] score_6_x42;
wire signed [DEBIT:0] score_6_x43;
wire signed [DEBIT:0] score_6_x44;
wire signed [DEBIT:0] score_6_x45;
wire signed [DEBIT:0] score_6_x46;
wire signed [DEBIT:0] score_6_x47;
wire signed [DEBIT:0] score_6_x48;
wire signed [DEBIT:0] score_6_x49;
wire signed [DEBIT:0] score_6_x50;
wire signed [DEBIT:0] score_6_x51;
wire signed [DEBIT:0] score_6_x52;
wire signed [DEBIT:0] score_6_x53;
wire signed [DEBIT:0] score_6_x54;
wire signed [DEBIT:0] score_6_x55;
wire signed [DEBIT:0] score_6_x56;
wire signed [DEBIT:0] score_6_x57;
wire signed [DEBIT:0] score_6_x58;
wire signed [DEBIT:0] score_6_x59;
wire signed [DEBIT:0] score_6_x60;
wire signed [DEBIT:0] score_6_x61;
wire signed [DEBIT:0] score_6_x62;
wire signed [DEBIT:0] score_6_x63;
wire signed [DEBIT:0] score_6_x64;
wire signed [DEBIT:0] score_6_x65;
wire signed [DEBIT:0] score_6_x66;
wire signed [DEBIT:0] score_6_x67;
wire signed [DEBIT:0] score_6_x68;
wire signed [DEBIT:0] score_6_x69;
wire signed [DEBIT:0] score_6_x70;
wire signed [DEBIT:0] score_6_x71;
wire signed [DEBIT:0] score_6_x72;
wire signed [DEBIT:0] score_6_x73;
wire signed [DEBIT:0] score_6_x74;
wire signed [DEBIT:0] score_6_x75;
wire signed [DEBIT:0] score_6_x76;
wire signed [DEBIT:0] score_6_x77;
wire signed [DEBIT:0] score_6_x78;
wire signed [DEBIT:0] score_6_x79;
wire signed [DEBIT:0] score_6_x80;
wire signed [DEBIT:0] score_6_x81;
wire signed [DEBIT:0] score_6_x82;
wire signed [DEBIT:0] score_6_x83;
wire signed [DEBIT:0] score_6_x84;
wire signed [DEBIT:0] score_6_x85;
wire signed [DEBIT:0] score_6_x86;
wire signed [DEBIT:0] score_6_x87;
wire signed [DEBIT:0] score_6_x88;
wire signed [DEBIT:0] score_6_x89;
wire signed [DEBIT:0] score_6_x90;
wire signed [DEBIT:0] score_6_x91;
wire signed [DEBIT:0] score_6_x92;
wire signed [DEBIT:0] score_6_x93;
wire signed [DEBIT:0] score_6_x94;
wire signed [DEBIT:0] score_6_x95;
wire signed [DEBIT:0] score_6_x96;
wire signed [DEBIT:0] score_6_x97;
wire signed [DEBIT:0] score_6_x98;
wire signed [DEBIT:0] score_6_x99;
wire signed [DEBIT:0] score_6_x100;
wire signed [DEBIT:0] score_6_x101;
wire signed [DEBIT:0] score_6_x102;
wire signed [DEBIT:0] score_6_x103;
wire signed [DEBIT:0] score_6_x104;
wire signed [DEBIT:0] score_6_x105;
wire signed [DEBIT:0] score_6_x106;
wire signed [DEBIT:0] score_6_x107;
wire signed [DEBIT:0] score_6_x108;
wire signed [DEBIT:0] score_6_x109;
wire signed [DEBIT:0] score_6_x110;
wire signed [DEBIT:0] score_6_x111;
wire signed [DEBIT:0] score_6_x112;
wire signed [DEBIT:0] score_6_x113;
wire signed [DEBIT:0] score_6_x114;
wire signed [DEBIT:0] score_6_x115;
wire signed [DEBIT:0] score_6_x116;
wire signed [DEBIT:0] score_6_x117;
wire signed [DEBIT:0] score_6_x118;
wire signed [DEBIT:0] score_6_x119;
wire signed [DEBIT:0] score_6_x120;
wire signed [DEBIT:0] score_6_x121;
wire signed [DEBIT:0] score_6_x122;
wire signed [DEBIT:0] score_6_x123;
wire signed [DEBIT:0] score_6_x124;
wire signed [DEBIT:0] score_6_x125;
wire signed [DEBIT:0] score_6_x126;
wire signed [DEBIT:0] score_6_x127;
wire signed [DEBIT:0] score_6_x128;
wire signed [DEBIT:0] score_6_x129;
wire signed [DEBIT:0] score_6_x130;
wire signed [DEBIT:0] score_6_x131;
wire signed [DEBIT:0] score_6_x132;
wire signed [DEBIT:0] score_6_x133;
wire signed [DEBIT:0] score_6_x134;
wire signed [DEBIT:0] score_6_x135;
wire signed [DEBIT:0] score_6_x136;
wire signed [DEBIT:0] score_6_x137;
wire signed [DEBIT:0] score_6_x138;
wire signed [DEBIT:0] score_6_x139;
wire signed [DEBIT:0] score_6_x140;
wire signed [DEBIT:0] score_6_x141;
wire signed [DEBIT:0] score_6_x142;
wire signed [DEBIT:0] score_6_x143;
wire signed [DEBIT:0] score_6_x144;
wire signed [DEBIT:0] score_6_x145;
wire signed [DEBIT:0] score_6_x146;
wire signed [DEBIT:0] score_6_x147;
wire signed [DEBIT:0] score_6_x148;
wire signed [DEBIT:0] score_6_x149;
wire signed [DEBIT:0] score_6_x150;
wire signed [DEBIT:0] score_6_x151;
wire signed [DEBIT:0] score_6_x152;
wire signed [DEBIT:0] score_6_x153;
wire signed [DEBIT:0] score_6_x154;
wire signed [DEBIT:0] score_6_x155;
wire signed [DEBIT:0] score_6_x156;
wire signed [DEBIT:0] score_6_x157;
wire signed [DEBIT:0] score_6_x158;
wire signed [DEBIT:0] score_6_x159;
wire signed [DEBIT:0] score_6_x160;
wire signed [DEBIT:0] score_6_x161;
wire signed [DEBIT:0] score_6_x162;
wire signed [DEBIT:0] score_6_x163;
wire signed [DEBIT:0] score_6_x164;
wire signed [DEBIT:0] score_6_x165;
wire signed [DEBIT:0] score_6_x166;
wire signed [DEBIT:0] score_6_x167;
wire signed [DEBIT:0] score_6_x168;
wire signed [DEBIT:0] score_6_x169;
wire signed [DEBIT:0] score_6_x170;
wire signed [DEBIT:0] score_6_x171;
wire signed [DEBIT:0] score_6_x172;
wire signed [DEBIT:0] score_6_x173;
wire signed [DEBIT:0] score_6_x174;
wire signed [DEBIT:0] score_6_x175;
wire signed [DEBIT:0] score_6_x176;
wire signed [DEBIT:0] score_6_x177;
wire signed [DEBIT:0] score_6_x178;
wire signed [DEBIT:0] score_6_x179;
wire signed [DEBIT:0] score_6_x180;
wire signed [DEBIT:0] score_6_x181;
wire signed [DEBIT:0] score_6_x182;
wire signed [DEBIT:0] score_6_x183;
wire signed [DEBIT:0] score_6_x184;
wire signed [DEBIT:0] score_6_x185;
wire signed [DEBIT:0] score_6_x186;
wire signed [DEBIT:0] score_6_x187;
wire signed [DEBIT:0] score_6_x188;
wire signed [DEBIT:0] score_6_x189;
wire signed [DEBIT:0] score_6_x190;
wire signed [DEBIT:0] score_6_x191;
wire signed [DEBIT:0] score_6_x192;
wire signed [DEBIT:0] score_6_x193;
wire signed [DEBIT:0] score_6_x194;
wire signed [DEBIT:0] score_6_x195;
wire signed [DEBIT:0] score_6_x196;
wire signed [DEBIT:0] score_6_x197;
wire signed [DEBIT:0] score_6_x198;
wire signed [DEBIT:0] score_6_x199;
wire signed [DEBIT:0] score_6_x200;
wire signed [DEBIT:0] score_6_x201;
wire signed [DEBIT:0] score_6_x202;
wire signed [DEBIT:0] score_6_x203;
wire signed [DEBIT:0] score_6_x204;
wire signed [DEBIT:0] score_6_x205;
wire signed [DEBIT:0] score_6_x206;
wire signed [DEBIT:0] score_6_x207;
wire signed [DEBIT:0] score_6_x208;
wire signed [DEBIT:0] score_6_x209;
wire signed [DEBIT:0] score_6_x210;
wire signed [DEBIT:0] score_6_x211;
wire signed [DEBIT:0] score_6_x212;
wire signed [DEBIT:0] score_6_x213;
wire signed [DEBIT:0] score_6_x214;
wire signed [DEBIT:0] score_6_x215;
wire signed [DEBIT:0] score_6_x216;
wire signed [DEBIT:0] score_6_x217;
wire signed [DEBIT:0] score_6_x218;
wire signed [DEBIT:0] score_6_x219;
wire signed [DEBIT:0] score_6_x220;
wire signed [DEBIT:0] score_6_x221;
wire signed [DEBIT:0] score_6_x222;
wire signed [DEBIT:0] score_6_x223;
wire signed [DEBIT:0] score_6_x224;
wire signed [DEBIT:0] score_6_x225;
wire signed [DEBIT:0] score_6_x226;
wire signed [DEBIT:0] score_6_x227;
wire signed [DEBIT:0] score_6_x228;
wire signed [DEBIT:0] score_6_x229;
wire signed [DEBIT:0] score_6_x230;
wire signed [DEBIT:0] score_6_x231;
wire signed [DEBIT:0] score_6_x232;
wire signed [DEBIT:0] score_6_x233;
wire signed [DEBIT:0] score_6_x234;
wire signed [DEBIT:0] score_6_x235;
wire signed [DEBIT:0] score_6_x236;
wire signed [DEBIT:0] score_6_x237;
wire signed [DEBIT:0] score_6_x238;
wire signed [DEBIT:0] score_6_x239;
wire signed [DEBIT:0] score_6_x240;
wire signed [DEBIT:0] score_6_x241;
wire signed [DEBIT:0] score_6_x242;
wire signed [DEBIT:0] score_6_x243;
wire signed [DEBIT:0] score_6_x244;
wire signed [DEBIT:0] score_6_x245;
wire signed [DEBIT:0] score_6_x246;
wire signed [DEBIT:0] score_6_x247;
wire signed [DEBIT:0] score_6_x248;
wire signed [DEBIT:0] score_6_x249;
wire signed [DEBIT:0] score_6_x250;
wire signed [DEBIT:0] score_6_x251;
wire signed [DEBIT:0] score_6_x252;
wire signed [DEBIT:0] score_6_x253;
wire signed [DEBIT:0] score_6_x254;
wire signed [DEBIT:0] score_6_x255;
wire signed [DEBIT:0] score_6_x256;
wire signed [DEBIT:0] score_6_x257;
wire signed [DEBIT:0] score_6_x258;
wire signed [DEBIT:0] score_6_x259;
wire signed [DEBIT:0] score_6_x260;
wire signed [DEBIT:0] score_6_x261;
wire signed [DEBIT:0] score_6_x262;
wire signed [DEBIT:0] score_6_x263;
wire signed [DEBIT:0] score_6_x264;
wire signed [DEBIT:0] score_6_x265;
wire signed [DEBIT:0] score_6_x266;
wire signed [DEBIT:0] score_6_x267;
wire signed [DEBIT:0] score_6_x268;
wire signed [DEBIT:0] score_6_x269;
wire signed [DEBIT:0] score_6_x270;
wire signed [DEBIT:0] score_6_x271;
wire signed [DEBIT:0] score_6_x272;
wire signed [DEBIT:0] score_6_x273;
wire signed [DEBIT:0] score_6_x274;
wire signed [DEBIT:0] score_6_x275;
wire signed [DEBIT:0] score_6_x276;
wire signed [DEBIT:0] score_6_x277;
wire signed [DEBIT:0] score_6_x278;
wire signed [DEBIT:0] score_6_x279;
wire signed [DEBIT:0] score_6_x280;
wire signed [DEBIT:0] score_6_x281;
wire signed [DEBIT:0] score_6_x282;
wire signed [DEBIT:0] score_6_x283;
wire signed [DEBIT:0] score_6_x284;
wire signed [DEBIT:0] score_6_x285;
wire signed [DEBIT:0] score_6_x286;
wire signed [DEBIT:0] score_6_x287;
wire signed [DEBIT:0] score_6_x288;
wire signed [DEBIT:0] score_6_x289;
wire signed [DEBIT:0] score_6_x290;
wire signed [DEBIT:0] score_6_x291;
wire signed [DEBIT:0] score_6_x292;
wire signed [DEBIT:0] score_6_x293;
wire signed [DEBIT:0] score_6_x294;
wire signed [DEBIT:0] score_6_x295;
wire signed [DEBIT:0] score_6_x296;
wire signed [DEBIT:0] score_6_x297;
wire signed [DEBIT:0] score_6_x298;
wire signed [DEBIT:0] score_6_x299;
wire signed [DEBIT:0] score_6_x300;
wire signed [DEBIT:0] score_6_x301;
wire signed [DEBIT:0] score_6_x302;
wire signed [DEBIT:0] score_6_x303;
wire signed [DEBIT:0] score_6_x304;
wire signed [DEBIT:0] score_6_x305;
wire signed [DEBIT:0] score_6_x306;
wire signed [DEBIT:0] score_6_x307;
wire signed [DEBIT:0] score_6_x308;
wire signed [DEBIT:0] score_6_x309;
wire signed [DEBIT:0] score_6_x310;
wire signed [DEBIT:0] score_6_x311;
wire signed [DEBIT:0] score_6_x312;
wire signed [DEBIT:0] score_6_x313;
wire signed [DEBIT:0] score_6_x314;
wire signed [DEBIT:0] score_6_x315;
wire signed [DEBIT:0] score_6_x316;
wire signed [DEBIT:0] score_6_x317;
wire signed [DEBIT:0] score_6_x318;
wire signed [DEBIT:0] score_6_x319;
wire signed [DEBIT:0] score_6_x320;
wire signed [DEBIT:0] score_6_x321;
wire signed [DEBIT:0] score_6_x322;
wire signed [DEBIT:0] score_6_x323;
wire signed [DEBIT:0] score_6_x324;
wire signed [DEBIT:0] score_6_x325;
wire signed [DEBIT:0] score_6_x326;
wire signed [DEBIT:0] score_6_x327;
wire signed [DEBIT:0] score_6_x328;
wire signed [DEBIT:0] score_6_x329;
wire signed [DEBIT:0] score_6_x330;
wire signed [DEBIT:0] score_6_x331;
wire signed [DEBIT:0] score_6_x332;
wire signed [DEBIT:0] score_6_x333;
wire signed [DEBIT:0] score_6_x334;
wire signed [DEBIT:0] score_6_x335;
wire signed [DEBIT:0] score_6_x336;
wire signed [DEBIT:0] score_6_x337;
wire signed [DEBIT:0] score_6_x338;
wire signed [DEBIT:0] score_6_x339;
wire signed [DEBIT:0] score_6_x340;
wire signed [DEBIT:0] score_6_x341;
wire signed [DEBIT:0] score_6_x342;
wire signed [DEBIT:0] score_6_x343;
wire signed [DEBIT:0] score_6_x344;
wire signed [DEBIT:0] score_6_x345;
wire signed [DEBIT:0] score_6_x346;
wire signed [DEBIT:0] score_6_x347;
wire signed [DEBIT:0] score_6_x348;
wire signed [DEBIT:0] score_6_x349;
wire signed [DEBIT:0] score_6_x350;
wire signed [DEBIT:0] score_6_x351;
wire signed [DEBIT:0] score_6_x352;
wire signed [DEBIT:0] score_6_x353;
wire signed [DEBIT:0] score_6_x354;
wire signed [DEBIT:0] score_6_x355;
wire signed [DEBIT:0] score_6_x356;
wire signed [DEBIT:0] score_6_x357;
wire signed [DEBIT:0] score_6_x358;
wire signed [DEBIT:0] score_6_x359;
wire signed [DEBIT:0] score_6_x360;
wire signed [DEBIT:0] score_6_x361;
wire signed [DEBIT:0] score_6_x362;
wire signed [DEBIT:0] score_6_x363;
wire signed [DEBIT:0] score_6_x364;
wire signed [DEBIT:0] score_6_x365;
wire signed [DEBIT:0] score_6_x366;
wire signed [DEBIT:0] score_6_x367;
wire signed [DEBIT:0] score_6_x368;
wire signed [DEBIT:0] score_6_x369;
wire signed [DEBIT:0] score_6_x370;
wire signed [DEBIT:0] score_6_x371;
wire signed [DEBIT:0] score_6_x372;
wire signed [DEBIT:0] score_6_x373;
wire signed [DEBIT:0] score_6_x374;
wire signed [DEBIT:0] score_6_x375;
wire signed [DEBIT:0] score_6_x376;
wire signed [DEBIT:0] score_6_x377;
wire signed [DEBIT:0] score_6_x378;
wire signed [DEBIT:0] score_6_x379;
wire signed [DEBIT:0] score_6_x380;
wire signed [DEBIT:0] score_6_x381;
wire signed [DEBIT:0] score_6_x382;
wire signed [DEBIT:0] score_6_x383;
wire signed [DEBIT:0] score_6_x384;
wire signed [DEBIT:0] score_6_x385;
wire signed [DEBIT:0] score_6_x386;
wire signed [DEBIT:0] score_6_x387;
wire signed [DEBIT:0] score_6_x388;
wire signed [DEBIT:0] score_6_x389;
wire signed [DEBIT:0] score_6_x390;
wire signed [DEBIT:0] score_6_x391;
wire signed [DEBIT:0] score_6_x392;
wire signed [DEBIT:0] score_6_x393;
wire signed [DEBIT:0] score_6_x394;
wire signed [DEBIT:0] score_6_x395;
wire signed [DEBIT:0] score_6_x396;
wire signed [DEBIT:0] score_6_x397;
wire signed [DEBIT:0] score_6_x398;
wire signed [DEBIT:0] score_6_x399;
wire signed [DEBIT:0] score_6_x400;
wire signed [DEBIT:0] score_6_x401;
wire signed [DEBIT:0] score_6_x402;
wire signed [DEBIT:0] score_6_x403;
wire signed [DEBIT:0] score_6_x404;
wire signed [DEBIT:0] score_6_x405;
wire signed [DEBIT:0] score_6_x406;
wire signed [DEBIT:0] score_6_x407;
wire signed [DEBIT:0] score_6_x408;
wire signed [DEBIT:0] score_6_x409;
wire signed [DEBIT:0] score_6_x410;
wire signed [DEBIT:0] score_6_x411;
wire signed [DEBIT:0] score_6_x412;
wire signed [DEBIT:0] score_6_x413;
wire signed [DEBIT:0] score_6_x414;
wire signed [DEBIT:0] score_6_x415;
wire signed [DEBIT:0] score_6_x416;
wire signed [DEBIT:0] score_6_x417;
wire signed [DEBIT:0] score_6_x418;
wire signed [DEBIT:0] score_6_x419;
wire signed [DEBIT:0] score_6_x420;
wire signed [DEBIT:0] score_6_x421;
wire signed [DEBIT:0] score_6_x422;
wire signed [DEBIT:0] score_6_x423;
wire signed [DEBIT:0] score_6_x424;
wire signed [DEBIT:0] score_6_x425;
wire signed [DEBIT:0] score_6_x426;
wire signed [DEBIT:0] score_6_x427;
wire signed [DEBIT:0] score_6_x428;
wire signed [DEBIT:0] score_6_x429;
wire signed [DEBIT:0] score_6_x430;
wire signed [DEBIT:0] score_6_x431;
wire signed [DEBIT:0] score_6_x432;
wire signed [DEBIT:0] score_6_x433;
wire signed [DEBIT:0] score_6_x434;
wire signed [DEBIT:0] score_6_x435;
wire signed [DEBIT:0] score_6_x436;
wire signed [DEBIT:0] score_6_x437;
wire signed [DEBIT:0] score_6_x438;
wire signed [DEBIT:0] score_6_x439;
wire signed [DEBIT:0] score_6_x440;
wire signed [DEBIT:0] score_6_x441;
wire signed [DEBIT:0] score_6_x442;
wire signed [DEBIT:0] score_6_x443;
wire signed [DEBIT:0] score_6_x444;
wire signed [DEBIT:0] score_6_x445;
wire signed [DEBIT:0] score_6_x446;
wire signed [DEBIT:0] score_6_x447;
wire signed [DEBIT:0] score_6_x448;
wire signed [DEBIT:0] score_6_x449;
wire signed [DEBIT:0] score_6_x450;
wire signed [DEBIT:0] score_6_x451;
wire signed [DEBIT:0] score_6_x452;
wire signed [DEBIT:0] score_6_x453;
wire signed [DEBIT:0] score_6_x454;
wire signed [DEBIT:0] score_6_x455;
wire signed [DEBIT:0] score_6_x456;
wire signed [DEBIT:0] score_6_x457;
wire signed [DEBIT:0] score_6_x458;
wire signed [DEBIT:0] score_6_x459;
wire signed [DEBIT:0] score_6_x460;
wire signed [DEBIT:0] score_6_x461;
wire signed [DEBIT:0] score_6_x462;
wire signed [DEBIT:0] score_6_x463;
wire signed [DEBIT:0] score_6_x464;
wire signed [DEBIT:0] score_6_x465;
wire signed [DEBIT:0] score_6_x466;
wire signed [DEBIT:0] score_6_x467;
wire signed [DEBIT:0] score_6_x468;
wire signed [DEBIT:0] score_6_x469;
wire signed [DEBIT:0] score_6_x470;
wire signed [DEBIT:0] score_6_x471;
wire signed [DEBIT:0] score_6_x472;
wire signed [DEBIT:0] score_6_x473;
wire signed [DEBIT:0] score_6_x474;
wire signed [DEBIT:0] score_6_x475;
wire signed [DEBIT:0] score_6_x476;
wire signed [DEBIT:0] score_6_x477;
wire signed [DEBIT:0] score_6_x478;
wire signed [DEBIT:0] score_6_x479;
wire signed [DEBIT:0] score_6_x480;
wire signed [DEBIT:0] score_6_x481;
wire signed [DEBIT:0] score_6_x482;
wire signed [DEBIT:0] score_6_x483;
wire signed [DEBIT:0] score_6_x484;
wire signed [DEBIT:0] score_6_x485;
wire signed [DEBIT:0] score_6_x486;
wire signed [DEBIT:0] score_6_x487;
wire signed [DEBIT:0] score_6_x488;
wire signed [DEBIT:0] score_6_x489;
wire signed [DEBIT:0] score_6_x490;
wire signed [DEBIT:0] score_6_x491;
wire signed [DEBIT:0] score_6_x492;
wire signed [DEBIT:0] score_6_x493;
wire signed [DEBIT:0] score_6_x494;
wire signed [DEBIT:0] score_6_x495;
wire signed [DEBIT:0] score_6_x496;
wire signed [DEBIT:0] score_6_x497;
wire signed [DEBIT:0] score_6_x498;
wire signed [DEBIT:0] score_6_x499;
wire signed [DEBIT:0] score_6_x500;
wire signed [DEBIT:0] score_6_x501;
wire signed [DEBIT:0] score_6_x502;
wire signed [DEBIT:0] score_6_x503;
wire signed [DEBIT:0] score_6_x504;
wire signed [DEBIT:0] score_6_x505;
wire signed [DEBIT:0] score_6_x506;
wire signed [DEBIT:0] score_6_x507;
wire signed [DEBIT:0] score_6_x508;
wire signed [DEBIT:0] score_6_x509;
wire signed [DEBIT:0] score_6_x510;
wire signed [DEBIT:0] score_6_x511;
wire signed [DEBIT:0] score_6_x512;
wire signed [DEBIT:0] score_6_x513;
wire signed [DEBIT:0] score_6_x514;
wire signed [DEBIT:0] score_6_x515;
wire signed [DEBIT:0] score_6_x516;
wire signed [DEBIT:0] score_6_x517;
wire signed [DEBIT:0] score_6_x518;
wire signed [DEBIT:0] score_6_x519;
wire signed [DEBIT:0] score_6_x520;
wire signed [DEBIT:0] score_6_x521;
wire signed [DEBIT:0] score_6_x522;
wire signed [DEBIT:0] score_6_x523;
wire signed [DEBIT:0] score_6_x524;
wire signed [DEBIT:0] score_6_x525;
wire signed [DEBIT:0] score_6_x526;
wire signed [DEBIT:0] score_6_x527;
wire signed [DEBIT:0] score_6_x528;
wire signed [DEBIT:0] score_6_x529;
wire signed [DEBIT:0] score_6_x530;
wire signed [DEBIT:0] score_6_x531;
wire signed [DEBIT:0] score_6_x532;
wire signed [DEBIT:0] score_6_x533;
wire signed [DEBIT:0] score_6_x534;
wire signed [DEBIT:0] score_6_x535;
wire signed [DEBIT:0] score_6_x536;
wire signed [DEBIT:0] score_6_x537;
wire signed [DEBIT:0] score_6_x538;
wire signed [DEBIT:0] score_6_x539;
wire signed [DEBIT:0] score_6_x540;
wire signed [DEBIT:0] score_6_x541;
wire signed [DEBIT:0] score_6_x542;
wire signed [DEBIT:0] score_6_x543;
wire signed [DEBIT:0] score_6_x544;
wire signed [DEBIT:0] score_6_x545;
wire signed [DEBIT:0] score_6_x546;
wire signed [DEBIT:0] score_6_x547;
wire signed [DEBIT:0] score_6_x548;
wire signed [DEBIT:0] score_6_x549;
wire signed [DEBIT:0] score_6_x550;
wire signed [DEBIT:0] score_6_x551;
wire signed [DEBIT:0] score_6_x552;
wire signed [DEBIT:0] score_6_x553;
wire signed [DEBIT:0] score_6_x554;
wire signed [DEBIT:0] score_6_x555;
wire signed [DEBIT:0] score_6_x556;
wire signed [DEBIT:0] score_6_x557;
wire signed [DEBIT:0] score_6_x558;
wire signed [DEBIT:0] score_6_x559;
wire signed [DEBIT:0] score_6_x560;
wire signed [DEBIT:0] score_6_x561;
wire signed [DEBIT:0] score_6_x562;
wire signed [DEBIT:0] score_6_x563;
wire signed [DEBIT:0] score_6_x564;
wire signed [DEBIT:0] score_6_x565;
wire signed [DEBIT:0] score_6_x566;
wire signed [DEBIT:0] score_6_x567;
wire signed [DEBIT:0] score_6_x568;
wire signed [DEBIT:0] score_6_x569;
wire signed [DEBIT:0] score_6_x570;
wire signed [DEBIT:0] score_6_x571;
wire signed [DEBIT:0] score_6_x572;
wire signed [DEBIT:0] score_6_x573;
wire signed [DEBIT:0] score_6_x574;
wire signed [DEBIT:0] score_6_x575;
wire signed [DEBIT:0] score_6_x576;
wire signed [DEBIT:0] score_6_x577;
wire signed [DEBIT:0] score_6_x578;
wire signed [DEBIT:0] score_6_x579;
wire signed [DEBIT:0] score_6_x580;
wire signed [DEBIT:0] score_6_x581;
wire signed [DEBIT:0] score_6_x582;
wire signed [DEBIT:0] score_6_x583;
wire signed [DEBIT:0] score_6_x584;
wire signed [DEBIT:0] score_6_x585;
wire signed [DEBIT:0] score_6_x586;
wire signed [DEBIT:0] score_6_x587;
wire signed [DEBIT:0] score_6_x588;
wire signed [DEBIT:0] score_6_x589;
wire signed [DEBIT:0] score_6_x590;
wire signed [DEBIT:0] score_6_x591;
wire signed [DEBIT:0] score_6_x592;
wire signed [DEBIT:0] score_6_x593;
wire signed [DEBIT:0] score_6_x594;
wire signed [DEBIT:0] score_6_x595;
wire signed [DEBIT:0] score_6_x596;
wire signed [DEBIT:0] score_6_x597;
wire signed [DEBIT:0] score_6_x598;
wire signed [DEBIT:0] score_6_x599;
wire signed [DEBIT:0] score_6_x600;
wire signed [DEBIT:0] score_6_x601;
wire signed [DEBIT:0] score_6_x602;
wire signed [DEBIT:0] score_6_x603;
wire signed [DEBIT:0] score_6_x604;
wire signed [DEBIT:0] score_6_x605;
wire signed [DEBIT:0] score_6_x606;
wire signed [DEBIT:0] score_6_x607;
wire signed [DEBIT:0] score_6_x608;
wire signed [DEBIT:0] score_6_x609;
wire signed [DEBIT:0] score_6_x610;
wire signed [DEBIT:0] score_6_x611;
wire signed [DEBIT:0] score_6_x612;
wire signed [DEBIT:0] score_6_x613;
wire signed [DEBIT:0] score_6_x614;
wire signed [DEBIT:0] score_6_x615;
wire signed [DEBIT:0] score_6_x616;
wire signed [DEBIT:0] score_6_x617;
wire signed [DEBIT:0] score_6_x618;
wire signed [DEBIT:0] score_6_x619;
wire signed [DEBIT:0] score_6_x620;
wire signed [DEBIT:0] score_6_x621;
wire signed [DEBIT:0] score_6_x622;
wire signed [DEBIT:0] score_6_x623;
wire signed [DEBIT:0] score_6_x624;
wire signed [DEBIT:0] score_6_x625;
wire signed [DEBIT:0] score_6_x626;
wire signed [DEBIT:0] score_6_x627;
wire signed [DEBIT:0] score_6_x628;
wire signed [DEBIT:0] score_6_x629;
wire signed [DEBIT:0] score_6_x630;
wire signed [DEBIT:0] score_6_x631;
wire signed [DEBIT:0] score_6_x632;
wire signed [DEBIT:0] score_6_x633;
wire signed [DEBIT:0] score_6_x634;
wire signed [DEBIT:0] score_6_x635;
wire signed [DEBIT:0] score_6_x636;
wire signed [DEBIT:0] score_6_x637;
wire signed [DEBIT:0] score_6_x638;
wire signed [DEBIT:0] score_6_x639;
wire signed [DEBIT:0] score_6_x640;
wire signed [DEBIT:0] score_6_x641;
wire signed [DEBIT:0] score_6_x642;
wire signed [DEBIT:0] score_6_x643;
wire signed [DEBIT:0] score_6_x644;
wire signed [DEBIT:0] score_6_x645;
wire signed [DEBIT:0] score_6_x646;
wire signed [DEBIT:0] score_6_x647;
wire signed [DEBIT:0] score_6_x648;
wire signed [DEBIT:0] score_6_x649;
wire signed [DEBIT:0] score_6_x650;
wire signed [DEBIT:0] score_6_x651;
wire signed [DEBIT:0] score_6_x652;
wire signed [DEBIT:0] score_6_x653;
wire signed [DEBIT:0] score_6_x654;
wire signed [DEBIT:0] score_6_x655;
wire signed [DEBIT:0] score_6_x656;
wire signed [DEBIT:0] score_6_x657;
wire signed [DEBIT:0] score_6_x658;
wire signed [DEBIT:0] score_6_x659;
wire signed [DEBIT:0] score_6_x660;
wire signed [DEBIT:0] score_6_x661;
wire signed [DEBIT:0] score_6_x662;
wire signed [DEBIT:0] score_6_x663;
wire signed [DEBIT:0] score_6_x664;
wire signed [DEBIT:0] score_6_x665;
wire signed [DEBIT:0] score_6_x666;
wire signed [DEBIT:0] score_6_x667;
wire signed [DEBIT:0] score_6_x668;
wire signed [DEBIT:0] score_6_x669;
wire signed [DEBIT:0] score_6_x670;
wire signed [DEBIT:0] score_6_x671;
wire signed [DEBIT:0] score_6_x672;
wire signed [DEBIT:0] score_6_x673;
wire signed [DEBIT:0] score_6_x674;
wire signed [DEBIT:0] score_6_x675;
wire signed [DEBIT:0] score_6_x676;
wire signed [DEBIT:0] score_6_x677;
wire signed [DEBIT:0] score_6_x678;
wire signed [DEBIT:0] score_6_x679;
wire signed [DEBIT:0] score_6_x680;
wire signed [DEBIT:0] score_6_x681;
wire signed [DEBIT:0] score_6_x682;
wire signed [DEBIT:0] score_6_x683;
wire signed [DEBIT:0] score_6_x684;
wire signed [DEBIT:0] score_6_x685;
wire signed [DEBIT:0] score_6_x686;
wire signed [DEBIT:0] score_6_x687;
wire signed [DEBIT:0] score_6_x688;
wire signed [DEBIT:0] score_6_x689;
wire signed [DEBIT:0] score_6_x690;
wire signed [DEBIT:0] score_6_x691;
wire signed [DEBIT:0] score_6_x692;
wire signed [DEBIT:0] score_6_x693;
wire signed [DEBIT:0] score_6_x694;
wire signed [DEBIT:0] score_6_x695;
wire signed [DEBIT:0] score_6_x696;
wire signed [DEBIT:0] score_6_x697;
wire signed [DEBIT:0] score_6_x698;
wire signed [DEBIT:0] score_6_x699;
wire signed [DEBIT:0] score_6_x700;
wire signed [DEBIT:0] score_6_x701;
wire signed [DEBIT:0] score_6_x702;
wire signed [DEBIT:0] score_6_x703;
wire signed [DEBIT:0] score_6_x704;
wire signed [DEBIT:0] score_6_x705;
wire signed [DEBIT:0] score_6_x706;
wire signed [DEBIT:0] score_6_x707;
wire signed [DEBIT:0] score_6_x708;
wire signed [DEBIT:0] score_6_x709;
wire signed [DEBIT:0] score_6_x710;
wire signed [DEBIT:0] score_6_x711;
wire signed [DEBIT:0] score_6_x712;
wire signed [DEBIT:0] score_6_x713;
wire signed [DEBIT:0] score_6_x714;
wire signed [DEBIT:0] score_6_x715;
wire signed [DEBIT:0] score_6_x716;
wire signed [DEBIT:0] score_6_x717;
wire signed [DEBIT:0] score_6_x718;
wire signed [DEBIT:0] score_6_x719;
wire signed [DEBIT:0] score_6_x720;
wire signed [DEBIT:0] score_6_x721;
wire signed [DEBIT:0] score_6_x722;
wire signed [DEBIT:0] score_6_x723;
wire signed [DEBIT:0] score_6_x724;
wire signed [DEBIT:0] score_6_x725;
wire signed [DEBIT:0] score_6_x726;
wire signed [DEBIT:0] score_6_x727;
wire signed [DEBIT:0] score_6_x728;
wire signed [DEBIT:0] score_6_x729;
wire signed [DEBIT:0] score_6_x730;
wire signed [DEBIT:0] score_6_x731;
wire signed [DEBIT:0] score_6_x732;
wire signed [DEBIT:0] score_6_x733;
wire signed [DEBIT:0] score_6_x734;
wire signed [DEBIT:0] score_6_x735;
wire signed [DEBIT:0] score_6_x736;
wire signed [DEBIT:0] score_6_x737;
wire signed [DEBIT:0] score_6_x738;
wire signed [DEBIT:0] score_6_x739;
wire signed [DEBIT:0] score_6_x740;
wire signed [DEBIT:0] score_6_x741;
wire signed [DEBIT:0] score_6_x742;
wire signed [DEBIT:0] score_6_x743;
wire signed [DEBIT:0] score_6_x744;
wire signed [DEBIT:0] score_6_x745;
wire signed [DEBIT:0] score_6_x746;
wire signed [DEBIT:0] score_6_x747;
wire signed [DEBIT:0] score_6_x748;
wire signed [DEBIT:0] score_6_x749;
wire signed [DEBIT:0] score_6_x750;
wire signed [DEBIT:0] score_6_x751;
wire signed [DEBIT:0] score_6_x752;
wire signed [DEBIT:0] score_6_x753;
wire signed [DEBIT:0] score_6_x754;
wire signed [DEBIT:0] score_6_x755;
wire signed [DEBIT:0] score_6_x756;
wire signed [DEBIT:0] score_6_x757;
wire signed [DEBIT:0] score_6_x758;
wire signed [DEBIT:0] score_6_x759;
wire signed [DEBIT:0] score_6_x760;
wire signed [DEBIT:0] score_6_x761;
wire signed [DEBIT:0] score_6_x762;
wire signed [DEBIT:0] score_6_x763;
wire signed [DEBIT:0] score_6_x764;
wire signed [DEBIT:0] score_6_x765;
wire signed [DEBIT:0] score_6_x766;
wire signed [DEBIT:0] score_6_x767;
wire signed [DEBIT:0] score_6_x768;
wire signed [DEBIT:0] score_6_x769;
wire signed [DEBIT:0] score_6_x770;
wire signed [DEBIT:0] score_6_x771;
wire signed [DEBIT:0] score_6_x772;
wire signed [DEBIT:0] score_6_x773;
wire signed [DEBIT:0] score_6_x774;
wire signed [DEBIT:0] score_6_x775;
wire signed [DEBIT:0] score_6_x776;
wire signed [DEBIT:0] score_6_x777;
wire signed [DEBIT:0] score_6_x778;
wire signed [DEBIT:0] score_6_x779;
wire signed [DEBIT:0] score_6_x780;
wire signed [DEBIT:0] score_6_x781;
wire signed [DEBIT:0] score_6_x782;
wire signed [DEBIT:0] score_6_x783;
wire signed [DEBIT:0] score_6_x784;
wire signed [DEBIT:0] score_7_x1;
wire signed [DEBIT:0] score_7_x2;
wire signed [DEBIT:0] score_7_x3;
wire signed [DEBIT:0] score_7_x4;
wire signed [DEBIT:0] score_7_x5;
wire signed [DEBIT:0] score_7_x6;
wire signed [DEBIT:0] score_7_x7;
wire signed [DEBIT:0] score_7_x8;
wire signed [DEBIT:0] score_7_x9;
wire signed [DEBIT:0] score_7_x10;
wire signed [DEBIT:0] score_7_x11;
wire signed [DEBIT:0] score_7_x12;
wire signed [DEBIT:0] score_7_x13;
wire signed [DEBIT:0] score_7_x14;
wire signed [DEBIT:0] score_7_x15;
wire signed [DEBIT:0] score_7_x16;
wire signed [DEBIT:0] score_7_x17;
wire signed [DEBIT:0] score_7_x18;
wire signed [DEBIT:0] score_7_x19;
wire signed [DEBIT:0] score_7_x20;
wire signed [DEBIT:0] score_7_x21;
wire signed [DEBIT:0] score_7_x22;
wire signed [DEBIT:0] score_7_x23;
wire signed [DEBIT:0] score_7_x24;
wire signed [DEBIT:0] score_7_x25;
wire signed [DEBIT:0] score_7_x26;
wire signed [DEBIT:0] score_7_x27;
wire signed [DEBIT:0] score_7_x28;
wire signed [DEBIT:0] score_7_x29;
wire signed [DEBIT:0] score_7_x30;
wire signed [DEBIT:0] score_7_x31;
wire signed [DEBIT:0] score_7_x32;
wire signed [DEBIT:0] score_7_x33;
wire signed [DEBIT:0] score_7_x34;
wire signed [DEBIT:0] score_7_x35;
wire signed [DEBIT:0] score_7_x36;
wire signed [DEBIT:0] score_7_x37;
wire signed [DEBIT:0] score_7_x38;
wire signed [DEBIT:0] score_7_x39;
wire signed [DEBIT:0] score_7_x40;
wire signed [DEBIT:0] score_7_x41;
wire signed [DEBIT:0] score_7_x42;
wire signed [DEBIT:0] score_7_x43;
wire signed [DEBIT:0] score_7_x44;
wire signed [DEBIT:0] score_7_x45;
wire signed [DEBIT:0] score_7_x46;
wire signed [DEBIT:0] score_7_x47;
wire signed [DEBIT:0] score_7_x48;
wire signed [DEBIT:0] score_7_x49;
wire signed [DEBIT:0] score_7_x50;
wire signed [DEBIT:0] score_7_x51;
wire signed [DEBIT:0] score_7_x52;
wire signed [DEBIT:0] score_7_x53;
wire signed [DEBIT:0] score_7_x54;
wire signed [DEBIT:0] score_7_x55;
wire signed [DEBIT:0] score_7_x56;
wire signed [DEBIT:0] score_7_x57;
wire signed [DEBIT:0] score_7_x58;
wire signed [DEBIT:0] score_7_x59;
wire signed [DEBIT:0] score_7_x60;
wire signed [DEBIT:0] score_7_x61;
wire signed [DEBIT:0] score_7_x62;
wire signed [DEBIT:0] score_7_x63;
wire signed [DEBIT:0] score_7_x64;
wire signed [DEBIT:0] score_7_x65;
wire signed [DEBIT:0] score_7_x66;
wire signed [DEBIT:0] score_7_x67;
wire signed [DEBIT:0] score_7_x68;
wire signed [DEBIT:0] score_7_x69;
wire signed [DEBIT:0] score_7_x70;
wire signed [DEBIT:0] score_7_x71;
wire signed [DEBIT:0] score_7_x72;
wire signed [DEBIT:0] score_7_x73;
wire signed [DEBIT:0] score_7_x74;
wire signed [DEBIT:0] score_7_x75;
wire signed [DEBIT:0] score_7_x76;
wire signed [DEBIT:0] score_7_x77;
wire signed [DEBIT:0] score_7_x78;
wire signed [DEBIT:0] score_7_x79;
wire signed [DEBIT:0] score_7_x80;
wire signed [DEBIT:0] score_7_x81;
wire signed [DEBIT:0] score_7_x82;
wire signed [DEBIT:0] score_7_x83;
wire signed [DEBIT:0] score_7_x84;
wire signed [DEBIT:0] score_7_x85;
wire signed [DEBIT:0] score_7_x86;
wire signed [DEBIT:0] score_7_x87;
wire signed [DEBIT:0] score_7_x88;
wire signed [DEBIT:0] score_7_x89;
wire signed [DEBIT:0] score_7_x90;
wire signed [DEBIT:0] score_7_x91;
wire signed [DEBIT:0] score_7_x92;
wire signed [DEBIT:0] score_7_x93;
wire signed [DEBIT:0] score_7_x94;
wire signed [DEBIT:0] score_7_x95;
wire signed [DEBIT:0] score_7_x96;
wire signed [DEBIT:0] score_7_x97;
wire signed [DEBIT:0] score_7_x98;
wire signed [DEBIT:0] score_7_x99;
wire signed [DEBIT:0] score_7_x100;
wire signed [DEBIT:0] score_7_x101;
wire signed [DEBIT:0] score_7_x102;
wire signed [DEBIT:0] score_7_x103;
wire signed [DEBIT:0] score_7_x104;
wire signed [DEBIT:0] score_7_x105;
wire signed [DEBIT:0] score_7_x106;
wire signed [DEBIT:0] score_7_x107;
wire signed [DEBIT:0] score_7_x108;
wire signed [DEBIT:0] score_7_x109;
wire signed [DEBIT:0] score_7_x110;
wire signed [DEBIT:0] score_7_x111;
wire signed [DEBIT:0] score_7_x112;
wire signed [DEBIT:0] score_7_x113;
wire signed [DEBIT:0] score_7_x114;
wire signed [DEBIT:0] score_7_x115;
wire signed [DEBIT:0] score_7_x116;
wire signed [DEBIT:0] score_7_x117;
wire signed [DEBIT:0] score_7_x118;
wire signed [DEBIT:0] score_7_x119;
wire signed [DEBIT:0] score_7_x120;
wire signed [DEBIT:0] score_7_x121;
wire signed [DEBIT:0] score_7_x122;
wire signed [DEBIT:0] score_7_x123;
wire signed [DEBIT:0] score_7_x124;
wire signed [DEBIT:0] score_7_x125;
wire signed [DEBIT:0] score_7_x126;
wire signed [DEBIT:0] score_7_x127;
wire signed [DEBIT:0] score_7_x128;
wire signed [DEBIT:0] score_7_x129;
wire signed [DEBIT:0] score_7_x130;
wire signed [DEBIT:0] score_7_x131;
wire signed [DEBIT:0] score_7_x132;
wire signed [DEBIT:0] score_7_x133;
wire signed [DEBIT:0] score_7_x134;
wire signed [DEBIT:0] score_7_x135;
wire signed [DEBIT:0] score_7_x136;
wire signed [DEBIT:0] score_7_x137;
wire signed [DEBIT:0] score_7_x138;
wire signed [DEBIT:0] score_7_x139;
wire signed [DEBIT:0] score_7_x140;
wire signed [DEBIT:0] score_7_x141;
wire signed [DEBIT:0] score_7_x142;
wire signed [DEBIT:0] score_7_x143;
wire signed [DEBIT:0] score_7_x144;
wire signed [DEBIT:0] score_7_x145;
wire signed [DEBIT:0] score_7_x146;
wire signed [DEBIT:0] score_7_x147;
wire signed [DEBIT:0] score_7_x148;
wire signed [DEBIT:0] score_7_x149;
wire signed [DEBIT:0] score_7_x150;
wire signed [DEBIT:0] score_7_x151;
wire signed [DEBIT:0] score_7_x152;
wire signed [DEBIT:0] score_7_x153;
wire signed [DEBIT:0] score_7_x154;
wire signed [DEBIT:0] score_7_x155;
wire signed [DEBIT:0] score_7_x156;
wire signed [DEBIT:0] score_7_x157;
wire signed [DEBIT:0] score_7_x158;
wire signed [DEBIT:0] score_7_x159;
wire signed [DEBIT:0] score_7_x160;
wire signed [DEBIT:0] score_7_x161;
wire signed [DEBIT:0] score_7_x162;
wire signed [DEBIT:0] score_7_x163;
wire signed [DEBIT:0] score_7_x164;
wire signed [DEBIT:0] score_7_x165;
wire signed [DEBIT:0] score_7_x166;
wire signed [DEBIT:0] score_7_x167;
wire signed [DEBIT:0] score_7_x168;
wire signed [DEBIT:0] score_7_x169;
wire signed [DEBIT:0] score_7_x170;
wire signed [DEBIT:0] score_7_x171;
wire signed [DEBIT:0] score_7_x172;
wire signed [DEBIT:0] score_7_x173;
wire signed [DEBIT:0] score_7_x174;
wire signed [DEBIT:0] score_7_x175;
wire signed [DEBIT:0] score_7_x176;
wire signed [DEBIT:0] score_7_x177;
wire signed [DEBIT:0] score_7_x178;
wire signed [DEBIT:0] score_7_x179;
wire signed [DEBIT:0] score_7_x180;
wire signed [DEBIT:0] score_7_x181;
wire signed [DEBIT:0] score_7_x182;
wire signed [DEBIT:0] score_7_x183;
wire signed [DEBIT:0] score_7_x184;
wire signed [DEBIT:0] score_7_x185;
wire signed [DEBIT:0] score_7_x186;
wire signed [DEBIT:0] score_7_x187;
wire signed [DEBIT:0] score_7_x188;
wire signed [DEBIT:0] score_7_x189;
wire signed [DEBIT:0] score_7_x190;
wire signed [DEBIT:0] score_7_x191;
wire signed [DEBIT:0] score_7_x192;
wire signed [DEBIT:0] score_7_x193;
wire signed [DEBIT:0] score_7_x194;
wire signed [DEBIT:0] score_7_x195;
wire signed [DEBIT:0] score_7_x196;
wire signed [DEBIT:0] score_7_x197;
wire signed [DEBIT:0] score_7_x198;
wire signed [DEBIT:0] score_7_x199;
wire signed [DEBIT:0] score_7_x200;
wire signed [DEBIT:0] score_7_x201;
wire signed [DEBIT:0] score_7_x202;
wire signed [DEBIT:0] score_7_x203;
wire signed [DEBIT:0] score_7_x204;
wire signed [DEBIT:0] score_7_x205;
wire signed [DEBIT:0] score_7_x206;
wire signed [DEBIT:0] score_7_x207;
wire signed [DEBIT:0] score_7_x208;
wire signed [DEBIT:0] score_7_x209;
wire signed [DEBIT:0] score_7_x210;
wire signed [DEBIT:0] score_7_x211;
wire signed [DEBIT:0] score_7_x212;
wire signed [DEBIT:0] score_7_x213;
wire signed [DEBIT:0] score_7_x214;
wire signed [DEBIT:0] score_7_x215;
wire signed [DEBIT:0] score_7_x216;
wire signed [DEBIT:0] score_7_x217;
wire signed [DEBIT:0] score_7_x218;
wire signed [DEBIT:0] score_7_x219;
wire signed [DEBIT:0] score_7_x220;
wire signed [DEBIT:0] score_7_x221;
wire signed [DEBIT:0] score_7_x222;
wire signed [DEBIT:0] score_7_x223;
wire signed [DEBIT:0] score_7_x224;
wire signed [DEBIT:0] score_7_x225;
wire signed [DEBIT:0] score_7_x226;
wire signed [DEBIT:0] score_7_x227;
wire signed [DEBIT:0] score_7_x228;
wire signed [DEBIT:0] score_7_x229;
wire signed [DEBIT:0] score_7_x230;
wire signed [DEBIT:0] score_7_x231;
wire signed [DEBIT:0] score_7_x232;
wire signed [DEBIT:0] score_7_x233;
wire signed [DEBIT:0] score_7_x234;
wire signed [DEBIT:0] score_7_x235;
wire signed [DEBIT:0] score_7_x236;
wire signed [DEBIT:0] score_7_x237;
wire signed [DEBIT:0] score_7_x238;
wire signed [DEBIT:0] score_7_x239;
wire signed [DEBIT:0] score_7_x240;
wire signed [DEBIT:0] score_7_x241;
wire signed [DEBIT:0] score_7_x242;
wire signed [DEBIT:0] score_7_x243;
wire signed [DEBIT:0] score_7_x244;
wire signed [DEBIT:0] score_7_x245;
wire signed [DEBIT:0] score_7_x246;
wire signed [DEBIT:0] score_7_x247;
wire signed [DEBIT:0] score_7_x248;
wire signed [DEBIT:0] score_7_x249;
wire signed [DEBIT:0] score_7_x250;
wire signed [DEBIT:0] score_7_x251;
wire signed [DEBIT:0] score_7_x252;
wire signed [DEBIT:0] score_7_x253;
wire signed [DEBIT:0] score_7_x254;
wire signed [DEBIT:0] score_7_x255;
wire signed [DEBIT:0] score_7_x256;
wire signed [DEBIT:0] score_7_x257;
wire signed [DEBIT:0] score_7_x258;
wire signed [DEBIT:0] score_7_x259;
wire signed [DEBIT:0] score_7_x260;
wire signed [DEBIT:0] score_7_x261;
wire signed [DEBIT:0] score_7_x262;
wire signed [DEBIT:0] score_7_x263;
wire signed [DEBIT:0] score_7_x264;
wire signed [DEBIT:0] score_7_x265;
wire signed [DEBIT:0] score_7_x266;
wire signed [DEBIT:0] score_7_x267;
wire signed [DEBIT:0] score_7_x268;
wire signed [DEBIT:0] score_7_x269;
wire signed [DEBIT:0] score_7_x270;
wire signed [DEBIT:0] score_7_x271;
wire signed [DEBIT:0] score_7_x272;
wire signed [DEBIT:0] score_7_x273;
wire signed [DEBIT:0] score_7_x274;
wire signed [DEBIT:0] score_7_x275;
wire signed [DEBIT:0] score_7_x276;
wire signed [DEBIT:0] score_7_x277;
wire signed [DEBIT:0] score_7_x278;
wire signed [DEBIT:0] score_7_x279;
wire signed [DEBIT:0] score_7_x280;
wire signed [DEBIT:0] score_7_x281;
wire signed [DEBIT:0] score_7_x282;
wire signed [DEBIT:0] score_7_x283;
wire signed [DEBIT:0] score_7_x284;
wire signed [DEBIT:0] score_7_x285;
wire signed [DEBIT:0] score_7_x286;
wire signed [DEBIT:0] score_7_x287;
wire signed [DEBIT:0] score_7_x288;
wire signed [DEBIT:0] score_7_x289;
wire signed [DEBIT:0] score_7_x290;
wire signed [DEBIT:0] score_7_x291;
wire signed [DEBIT:0] score_7_x292;
wire signed [DEBIT:0] score_7_x293;
wire signed [DEBIT:0] score_7_x294;
wire signed [DEBIT:0] score_7_x295;
wire signed [DEBIT:0] score_7_x296;
wire signed [DEBIT:0] score_7_x297;
wire signed [DEBIT:0] score_7_x298;
wire signed [DEBIT:0] score_7_x299;
wire signed [DEBIT:0] score_7_x300;
wire signed [DEBIT:0] score_7_x301;
wire signed [DEBIT:0] score_7_x302;
wire signed [DEBIT:0] score_7_x303;
wire signed [DEBIT:0] score_7_x304;
wire signed [DEBIT:0] score_7_x305;
wire signed [DEBIT:0] score_7_x306;
wire signed [DEBIT:0] score_7_x307;
wire signed [DEBIT:0] score_7_x308;
wire signed [DEBIT:0] score_7_x309;
wire signed [DEBIT:0] score_7_x310;
wire signed [DEBIT:0] score_7_x311;
wire signed [DEBIT:0] score_7_x312;
wire signed [DEBIT:0] score_7_x313;
wire signed [DEBIT:0] score_7_x314;
wire signed [DEBIT:0] score_7_x315;
wire signed [DEBIT:0] score_7_x316;
wire signed [DEBIT:0] score_7_x317;
wire signed [DEBIT:0] score_7_x318;
wire signed [DEBIT:0] score_7_x319;
wire signed [DEBIT:0] score_7_x320;
wire signed [DEBIT:0] score_7_x321;
wire signed [DEBIT:0] score_7_x322;
wire signed [DEBIT:0] score_7_x323;
wire signed [DEBIT:0] score_7_x324;
wire signed [DEBIT:0] score_7_x325;
wire signed [DEBIT:0] score_7_x326;
wire signed [DEBIT:0] score_7_x327;
wire signed [DEBIT:0] score_7_x328;
wire signed [DEBIT:0] score_7_x329;
wire signed [DEBIT:0] score_7_x330;
wire signed [DEBIT:0] score_7_x331;
wire signed [DEBIT:0] score_7_x332;
wire signed [DEBIT:0] score_7_x333;
wire signed [DEBIT:0] score_7_x334;
wire signed [DEBIT:0] score_7_x335;
wire signed [DEBIT:0] score_7_x336;
wire signed [DEBIT:0] score_7_x337;
wire signed [DEBIT:0] score_7_x338;
wire signed [DEBIT:0] score_7_x339;
wire signed [DEBIT:0] score_7_x340;
wire signed [DEBIT:0] score_7_x341;
wire signed [DEBIT:0] score_7_x342;
wire signed [DEBIT:0] score_7_x343;
wire signed [DEBIT:0] score_7_x344;
wire signed [DEBIT:0] score_7_x345;
wire signed [DEBIT:0] score_7_x346;
wire signed [DEBIT:0] score_7_x347;
wire signed [DEBIT:0] score_7_x348;
wire signed [DEBIT:0] score_7_x349;
wire signed [DEBIT:0] score_7_x350;
wire signed [DEBIT:0] score_7_x351;
wire signed [DEBIT:0] score_7_x352;
wire signed [DEBIT:0] score_7_x353;
wire signed [DEBIT:0] score_7_x354;
wire signed [DEBIT:0] score_7_x355;
wire signed [DEBIT:0] score_7_x356;
wire signed [DEBIT:0] score_7_x357;
wire signed [DEBIT:0] score_7_x358;
wire signed [DEBIT:0] score_7_x359;
wire signed [DEBIT:0] score_7_x360;
wire signed [DEBIT:0] score_7_x361;
wire signed [DEBIT:0] score_7_x362;
wire signed [DEBIT:0] score_7_x363;
wire signed [DEBIT:0] score_7_x364;
wire signed [DEBIT:0] score_7_x365;
wire signed [DEBIT:0] score_7_x366;
wire signed [DEBIT:0] score_7_x367;
wire signed [DEBIT:0] score_7_x368;
wire signed [DEBIT:0] score_7_x369;
wire signed [DEBIT:0] score_7_x370;
wire signed [DEBIT:0] score_7_x371;
wire signed [DEBIT:0] score_7_x372;
wire signed [DEBIT:0] score_7_x373;
wire signed [DEBIT:0] score_7_x374;
wire signed [DEBIT:0] score_7_x375;
wire signed [DEBIT:0] score_7_x376;
wire signed [DEBIT:0] score_7_x377;
wire signed [DEBIT:0] score_7_x378;
wire signed [DEBIT:0] score_7_x379;
wire signed [DEBIT:0] score_7_x380;
wire signed [DEBIT:0] score_7_x381;
wire signed [DEBIT:0] score_7_x382;
wire signed [DEBIT:0] score_7_x383;
wire signed [DEBIT:0] score_7_x384;
wire signed [DEBIT:0] score_7_x385;
wire signed [DEBIT:0] score_7_x386;
wire signed [DEBIT:0] score_7_x387;
wire signed [DEBIT:0] score_7_x388;
wire signed [DEBIT:0] score_7_x389;
wire signed [DEBIT:0] score_7_x390;
wire signed [DEBIT:0] score_7_x391;
wire signed [DEBIT:0] score_7_x392;
wire signed [DEBIT:0] score_7_x393;
wire signed [DEBIT:0] score_7_x394;
wire signed [DEBIT:0] score_7_x395;
wire signed [DEBIT:0] score_7_x396;
wire signed [DEBIT:0] score_7_x397;
wire signed [DEBIT:0] score_7_x398;
wire signed [DEBIT:0] score_7_x399;
wire signed [DEBIT:0] score_7_x400;
wire signed [DEBIT:0] score_7_x401;
wire signed [DEBIT:0] score_7_x402;
wire signed [DEBIT:0] score_7_x403;
wire signed [DEBIT:0] score_7_x404;
wire signed [DEBIT:0] score_7_x405;
wire signed [DEBIT:0] score_7_x406;
wire signed [DEBIT:0] score_7_x407;
wire signed [DEBIT:0] score_7_x408;
wire signed [DEBIT:0] score_7_x409;
wire signed [DEBIT:0] score_7_x410;
wire signed [DEBIT:0] score_7_x411;
wire signed [DEBIT:0] score_7_x412;
wire signed [DEBIT:0] score_7_x413;
wire signed [DEBIT:0] score_7_x414;
wire signed [DEBIT:0] score_7_x415;
wire signed [DEBIT:0] score_7_x416;
wire signed [DEBIT:0] score_7_x417;
wire signed [DEBIT:0] score_7_x418;
wire signed [DEBIT:0] score_7_x419;
wire signed [DEBIT:0] score_7_x420;
wire signed [DEBIT:0] score_7_x421;
wire signed [DEBIT:0] score_7_x422;
wire signed [DEBIT:0] score_7_x423;
wire signed [DEBIT:0] score_7_x424;
wire signed [DEBIT:0] score_7_x425;
wire signed [DEBIT:0] score_7_x426;
wire signed [DEBIT:0] score_7_x427;
wire signed [DEBIT:0] score_7_x428;
wire signed [DEBIT:0] score_7_x429;
wire signed [DEBIT:0] score_7_x430;
wire signed [DEBIT:0] score_7_x431;
wire signed [DEBIT:0] score_7_x432;
wire signed [DEBIT:0] score_7_x433;
wire signed [DEBIT:0] score_7_x434;
wire signed [DEBIT:0] score_7_x435;
wire signed [DEBIT:0] score_7_x436;
wire signed [DEBIT:0] score_7_x437;
wire signed [DEBIT:0] score_7_x438;
wire signed [DEBIT:0] score_7_x439;
wire signed [DEBIT:0] score_7_x440;
wire signed [DEBIT:0] score_7_x441;
wire signed [DEBIT:0] score_7_x442;
wire signed [DEBIT:0] score_7_x443;
wire signed [DEBIT:0] score_7_x444;
wire signed [DEBIT:0] score_7_x445;
wire signed [DEBIT:0] score_7_x446;
wire signed [DEBIT:0] score_7_x447;
wire signed [DEBIT:0] score_7_x448;
wire signed [DEBIT:0] score_7_x449;
wire signed [DEBIT:0] score_7_x450;
wire signed [DEBIT:0] score_7_x451;
wire signed [DEBIT:0] score_7_x452;
wire signed [DEBIT:0] score_7_x453;
wire signed [DEBIT:0] score_7_x454;
wire signed [DEBIT:0] score_7_x455;
wire signed [DEBIT:0] score_7_x456;
wire signed [DEBIT:0] score_7_x457;
wire signed [DEBIT:0] score_7_x458;
wire signed [DEBIT:0] score_7_x459;
wire signed [DEBIT:0] score_7_x460;
wire signed [DEBIT:0] score_7_x461;
wire signed [DEBIT:0] score_7_x462;
wire signed [DEBIT:0] score_7_x463;
wire signed [DEBIT:0] score_7_x464;
wire signed [DEBIT:0] score_7_x465;
wire signed [DEBIT:0] score_7_x466;
wire signed [DEBIT:0] score_7_x467;
wire signed [DEBIT:0] score_7_x468;
wire signed [DEBIT:0] score_7_x469;
wire signed [DEBIT:0] score_7_x470;
wire signed [DEBIT:0] score_7_x471;
wire signed [DEBIT:0] score_7_x472;
wire signed [DEBIT:0] score_7_x473;
wire signed [DEBIT:0] score_7_x474;
wire signed [DEBIT:0] score_7_x475;
wire signed [DEBIT:0] score_7_x476;
wire signed [DEBIT:0] score_7_x477;
wire signed [DEBIT:0] score_7_x478;
wire signed [DEBIT:0] score_7_x479;
wire signed [DEBIT:0] score_7_x480;
wire signed [DEBIT:0] score_7_x481;
wire signed [DEBIT:0] score_7_x482;
wire signed [DEBIT:0] score_7_x483;
wire signed [DEBIT:0] score_7_x484;
wire signed [DEBIT:0] score_7_x485;
wire signed [DEBIT:0] score_7_x486;
wire signed [DEBIT:0] score_7_x487;
wire signed [DEBIT:0] score_7_x488;
wire signed [DEBIT:0] score_7_x489;
wire signed [DEBIT:0] score_7_x490;
wire signed [DEBIT:0] score_7_x491;
wire signed [DEBIT:0] score_7_x492;
wire signed [DEBIT:0] score_7_x493;
wire signed [DEBIT:0] score_7_x494;
wire signed [DEBIT:0] score_7_x495;
wire signed [DEBIT:0] score_7_x496;
wire signed [DEBIT:0] score_7_x497;
wire signed [DEBIT:0] score_7_x498;
wire signed [DEBIT:0] score_7_x499;
wire signed [DEBIT:0] score_7_x500;
wire signed [DEBIT:0] score_7_x501;
wire signed [DEBIT:0] score_7_x502;
wire signed [DEBIT:0] score_7_x503;
wire signed [DEBIT:0] score_7_x504;
wire signed [DEBIT:0] score_7_x505;
wire signed [DEBIT:0] score_7_x506;
wire signed [DEBIT:0] score_7_x507;
wire signed [DEBIT:0] score_7_x508;
wire signed [DEBIT:0] score_7_x509;
wire signed [DEBIT:0] score_7_x510;
wire signed [DEBIT:0] score_7_x511;
wire signed [DEBIT:0] score_7_x512;
wire signed [DEBIT:0] score_7_x513;
wire signed [DEBIT:0] score_7_x514;
wire signed [DEBIT:0] score_7_x515;
wire signed [DEBIT:0] score_7_x516;
wire signed [DEBIT:0] score_7_x517;
wire signed [DEBIT:0] score_7_x518;
wire signed [DEBIT:0] score_7_x519;
wire signed [DEBIT:0] score_7_x520;
wire signed [DEBIT:0] score_7_x521;
wire signed [DEBIT:0] score_7_x522;
wire signed [DEBIT:0] score_7_x523;
wire signed [DEBIT:0] score_7_x524;
wire signed [DEBIT:0] score_7_x525;
wire signed [DEBIT:0] score_7_x526;
wire signed [DEBIT:0] score_7_x527;
wire signed [DEBIT:0] score_7_x528;
wire signed [DEBIT:0] score_7_x529;
wire signed [DEBIT:0] score_7_x530;
wire signed [DEBIT:0] score_7_x531;
wire signed [DEBIT:0] score_7_x532;
wire signed [DEBIT:0] score_7_x533;
wire signed [DEBIT:0] score_7_x534;
wire signed [DEBIT:0] score_7_x535;
wire signed [DEBIT:0] score_7_x536;
wire signed [DEBIT:0] score_7_x537;
wire signed [DEBIT:0] score_7_x538;
wire signed [DEBIT:0] score_7_x539;
wire signed [DEBIT:0] score_7_x540;
wire signed [DEBIT:0] score_7_x541;
wire signed [DEBIT:0] score_7_x542;
wire signed [DEBIT:0] score_7_x543;
wire signed [DEBIT:0] score_7_x544;
wire signed [DEBIT:0] score_7_x545;
wire signed [DEBIT:0] score_7_x546;
wire signed [DEBIT:0] score_7_x547;
wire signed [DEBIT:0] score_7_x548;
wire signed [DEBIT:0] score_7_x549;
wire signed [DEBIT:0] score_7_x550;
wire signed [DEBIT:0] score_7_x551;
wire signed [DEBIT:0] score_7_x552;
wire signed [DEBIT:0] score_7_x553;
wire signed [DEBIT:0] score_7_x554;
wire signed [DEBIT:0] score_7_x555;
wire signed [DEBIT:0] score_7_x556;
wire signed [DEBIT:0] score_7_x557;
wire signed [DEBIT:0] score_7_x558;
wire signed [DEBIT:0] score_7_x559;
wire signed [DEBIT:0] score_7_x560;
wire signed [DEBIT:0] score_7_x561;
wire signed [DEBIT:0] score_7_x562;
wire signed [DEBIT:0] score_7_x563;
wire signed [DEBIT:0] score_7_x564;
wire signed [DEBIT:0] score_7_x565;
wire signed [DEBIT:0] score_7_x566;
wire signed [DEBIT:0] score_7_x567;
wire signed [DEBIT:0] score_7_x568;
wire signed [DEBIT:0] score_7_x569;
wire signed [DEBIT:0] score_7_x570;
wire signed [DEBIT:0] score_7_x571;
wire signed [DEBIT:0] score_7_x572;
wire signed [DEBIT:0] score_7_x573;
wire signed [DEBIT:0] score_7_x574;
wire signed [DEBIT:0] score_7_x575;
wire signed [DEBIT:0] score_7_x576;
wire signed [DEBIT:0] score_7_x577;
wire signed [DEBIT:0] score_7_x578;
wire signed [DEBIT:0] score_7_x579;
wire signed [DEBIT:0] score_7_x580;
wire signed [DEBIT:0] score_7_x581;
wire signed [DEBIT:0] score_7_x582;
wire signed [DEBIT:0] score_7_x583;
wire signed [DEBIT:0] score_7_x584;
wire signed [DEBIT:0] score_7_x585;
wire signed [DEBIT:0] score_7_x586;
wire signed [DEBIT:0] score_7_x587;
wire signed [DEBIT:0] score_7_x588;
wire signed [DEBIT:0] score_7_x589;
wire signed [DEBIT:0] score_7_x590;
wire signed [DEBIT:0] score_7_x591;
wire signed [DEBIT:0] score_7_x592;
wire signed [DEBIT:0] score_7_x593;
wire signed [DEBIT:0] score_7_x594;
wire signed [DEBIT:0] score_7_x595;
wire signed [DEBIT:0] score_7_x596;
wire signed [DEBIT:0] score_7_x597;
wire signed [DEBIT:0] score_7_x598;
wire signed [DEBIT:0] score_7_x599;
wire signed [DEBIT:0] score_7_x600;
wire signed [DEBIT:0] score_7_x601;
wire signed [DEBIT:0] score_7_x602;
wire signed [DEBIT:0] score_7_x603;
wire signed [DEBIT:0] score_7_x604;
wire signed [DEBIT:0] score_7_x605;
wire signed [DEBIT:0] score_7_x606;
wire signed [DEBIT:0] score_7_x607;
wire signed [DEBIT:0] score_7_x608;
wire signed [DEBIT:0] score_7_x609;
wire signed [DEBIT:0] score_7_x610;
wire signed [DEBIT:0] score_7_x611;
wire signed [DEBIT:0] score_7_x612;
wire signed [DEBIT:0] score_7_x613;
wire signed [DEBIT:0] score_7_x614;
wire signed [DEBIT:0] score_7_x615;
wire signed [DEBIT:0] score_7_x616;
wire signed [DEBIT:0] score_7_x617;
wire signed [DEBIT:0] score_7_x618;
wire signed [DEBIT:0] score_7_x619;
wire signed [DEBIT:0] score_7_x620;
wire signed [DEBIT:0] score_7_x621;
wire signed [DEBIT:0] score_7_x622;
wire signed [DEBIT:0] score_7_x623;
wire signed [DEBIT:0] score_7_x624;
wire signed [DEBIT:0] score_7_x625;
wire signed [DEBIT:0] score_7_x626;
wire signed [DEBIT:0] score_7_x627;
wire signed [DEBIT:0] score_7_x628;
wire signed [DEBIT:0] score_7_x629;
wire signed [DEBIT:0] score_7_x630;
wire signed [DEBIT:0] score_7_x631;
wire signed [DEBIT:0] score_7_x632;
wire signed [DEBIT:0] score_7_x633;
wire signed [DEBIT:0] score_7_x634;
wire signed [DEBIT:0] score_7_x635;
wire signed [DEBIT:0] score_7_x636;
wire signed [DEBIT:0] score_7_x637;
wire signed [DEBIT:0] score_7_x638;
wire signed [DEBIT:0] score_7_x639;
wire signed [DEBIT:0] score_7_x640;
wire signed [DEBIT:0] score_7_x641;
wire signed [DEBIT:0] score_7_x642;
wire signed [DEBIT:0] score_7_x643;
wire signed [DEBIT:0] score_7_x644;
wire signed [DEBIT:0] score_7_x645;
wire signed [DEBIT:0] score_7_x646;
wire signed [DEBIT:0] score_7_x647;
wire signed [DEBIT:0] score_7_x648;
wire signed [DEBIT:0] score_7_x649;
wire signed [DEBIT:0] score_7_x650;
wire signed [DEBIT:0] score_7_x651;
wire signed [DEBIT:0] score_7_x652;
wire signed [DEBIT:0] score_7_x653;
wire signed [DEBIT:0] score_7_x654;
wire signed [DEBIT:0] score_7_x655;
wire signed [DEBIT:0] score_7_x656;
wire signed [DEBIT:0] score_7_x657;
wire signed [DEBIT:0] score_7_x658;
wire signed [DEBIT:0] score_7_x659;
wire signed [DEBIT:0] score_7_x660;
wire signed [DEBIT:0] score_7_x661;
wire signed [DEBIT:0] score_7_x662;
wire signed [DEBIT:0] score_7_x663;
wire signed [DEBIT:0] score_7_x664;
wire signed [DEBIT:0] score_7_x665;
wire signed [DEBIT:0] score_7_x666;
wire signed [DEBIT:0] score_7_x667;
wire signed [DEBIT:0] score_7_x668;
wire signed [DEBIT:0] score_7_x669;
wire signed [DEBIT:0] score_7_x670;
wire signed [DEBIT:0] score_7_x671;
wire signed [DEBIT:0] score_7_x672;
wire signed [DEBIT:0] score_7_x673;
wire signed [DEBIT:0] score_7_x674;
wire signed [DEBIT:0] score_7_x675;
wire signed [DEBIT:0] score_7_x676;
wire signed [DEBIT:0] score_7_x677;
wire signed [DEBIT:0] score_7_x678;
wire signed [DEBIT:0] score_7_x679;
wire signed [DEBIT:0] score_7_x680;
wire signed [DEBIT:0] score_7_x681;
wire signed [DEBIT:0] score_7_x682;
wire signed [DEBIT:0] score_7_x683;
wire signed [DEBIT:0] score_7_x684;
wire signed [DEBIT:0] score_7_x685;
wire signed [DEBIT:0] score_7_x686;
wire signed [DEBIT:0] score_7_x687;
wire signed [DEBIT:0] score_7_x688;
wire signed [DEBIT:0] score_7_x689;
wire signed [DEBIT:0] score_7_x690;
wire signed [DEBIT:0] score_7_x691;
wire signed [DEBIT:0] score_7_x692;
wire signed [DEBIT:0] score_7_x693;
wire signed [DEBIT:0] score_7_x694;
wire signed [DEBIT:0] score_7_x695;
wire signed [DEBIT:0] score_7_x696;
wire signed [DEBIT:0] score_7_x697;
wire signed [DEBIT:0] score_7_x698;
wire signed [DEBIT:0] score_7_x699;
wire signed [DEBIT:0] score_7_x700;
wire signed [DEBIT:0] score_7_x701;
wire signed [DEBIT:0] score_7_x702;
wire signed [DEBIT:0] score_7_x703;
wire signed [DEBIT:0] score_7_x704;
wire signed [DEBIT:0] score_7_x705;
wire signed [DEBIT:0] score_7_x706;
wire signed [DEBIT:0] score_7_x707;
wire signed [DEBIT:0] score_7_x708;
wire signed [DEBIT:0] score_7_x709;
wire signed [DEBIT:0] score_7_x710;
wire signed [DEBIT:0] score_7_x711;
wire signed [DEBIT:0] score_7_x712;
wire signed [DEBIT:0] score_7_x713;
wire signed [DEBIT:0] score_7_x714;
wire signed [DEBIT:0] score_7_x715;
wire signed [DEBIT:0] score_7_x716;
wire signed [DEBIT:0] score_7_x717;
wire signed [DEBIT:0] score_7_x718;
wire signed [DEBIT:0] score_7_x719;
wire signed [DEBIT:0] score_7_x720;
wire signed [DEBIT:0] score_7_x721;
wire signed [DEBIT:0] score_7_x722;
wire signed [DEBIT:0] score_7_x723;
wire signed [DEBIT:0] score_7_x724;
wire signed [DEBIT:0] score_7_x725;
wire signed [DEBIT:0] score_7_x726;
wire signed [DEBIT:0] score_7_x727;
wire signed [DEBIT:0] score_7_x728;
wire signed [DEBIT:0] score_7_x729;
wire signed [DEBIT:0] score_7_x730;
wire signed [DEBIT:0] score_7_x731;
wire signed [DEBIT:0] score_7_x732;
wire signed [DEBIT:0] score_7_x733;
wire signed [DEBIT:0] score_7_x734;
wire signed [DEBIT:0] score_7_x735;
wire signed [DEBIT:0] score_7_x736;
wire signed [DEBIT:0] score_7_x737;
wire signed [DEBIT:0] score_7_x738;
wire signed [DEBIT:0] score_7_x739;
wire signed [DEBIT:0] score_7_x740;
wire signed [DEBIT:0] score_7_x741;
wire signed [DEBIT:0] score_7_x742;
wire signed [DEBIT:0] score_7_x743;
wire signed [DEBIT:0] score_7_x744;
wire signed [DEBIT:0] score_7_x745;
wire signed [DEBIT:0] score_7_x746;
wire signed [DEBIT:0] score_7_x747;
wire signed [DEBIT:0] score_7_x748;
wire signed [DEBIT:0] score_7_x749;
wire signed [DEBIT:0] score_7_x750;
wire signed [DEBIT:0] score_7_x751;
wire signed [DEBIT:0] score_7_x752;
wire signed [DEBIT:0] score_7_x753;
wire signed [DEBIT:0] score_7_x754;
wire signed [DEBIT:0] score_7_x755;
wire signed [DEBIT:0] score_7_x756;
wire signed [DEBIT:0] score_7_x757;
wire signed [DEBIT:0] score_7_x758;
wire signed [DEBIT:0] score_7_x759;
wire signed [DEBIT:0] score_7_x760;
wire signed [DEBIT:0] score_7_x761;
wire signed [DEBIT:0] score_7_x762;
wire signed [DEBIT:0] score_7_x763;
wire signed [DEBIT:0] score_7_x764;
wire signed [DEBIT:0] score_7_x765;
wire signed [DEBIT:0] score_7_x766;
wire signed [DEBIT:0] score_7_x767;
wire signed [DEBIT:0] score_7_x768;
wire signed [DEBIT:0] score_7_x769;
wire signed [DEBIT:0] score_7_x770;
wire signed [DEBIT:0] score_7_x771;
wire signed [DEBIT:0] score_7_x772;
wire signed [DEBIT:0] score_7_x773;
wire signed [DEBIT:0] score_7_x774;
wire signed [DEBIT:0] score_7_x775;
wire signed [DEBIT:0] score_7_x776;
wire signed [DEBIT:0] score_7_x777;
wire signed [DEBIT:0] score_7_x778;
wire signed [DEBIT:0] score_7_x779;
wire signed [DEBIT:0] score_7_x780;
wire signed [DEBIT:0] score_7_x781;
wire signed [DEBIT:0] score_7_x782;
wire signed [DEBIT:0] score_7_x783;
wire signed [DEBIT:0] score_7_x784;
wire signed [DEBIT:0] score_8_x1;
wire signed [DEBIT:0] score_8_x2;
wire signed [DEBIT:0] score_8_x3;
wire signed [DEBIT:0] score_8_x4;
wire signed [DEBIT:0] score_8_x5;
wire signed [DEBIT:0] score_8_x6;
wire signed [DEBIT:0] score_8_x7;
wire signed [DEBIT:0] score_8_x8;
wire signed [DEBIT:0] score_8_x9;
wire signed [DEBIT:0] score_8_x10;
wire signed [DEBIT:0] score_8_x11;
wire signed [DEBIT:0] score_8_x12;
wire signed [DEBIT:0] score_8_x13;
wire signed [DEBIT:0] score_8_x14;
wire signed [DEBIT:0] score_8_x15;
wire signed [DEBIT:0] score_8_x16;
wire signed [DEBIT:0] score_8_x17;
wire signed [DEBIT:0] score_8_x18;
wire signed [DEBIT:0] score_8_x19;
wire signed [DEBIT:0] score_8_x20;
wire signed [DEBIT:0] score_8_x21;
wire signed [DEBIT:0] score_8_x22;
wire signed [DEBIT:0] score_8_x23;
wire signed [DEBIT:0] score_8_x24;
wire signed [DEBIT:0] score_8_x25;
wire signed [DEBIT:0] score_8_x26;
wire signed [DEBIT:0] score_8_x27;
wire signed [DEBIT:0] score_8_x28;
wire signed [DEBIT:0] score_8_x29;
wire signed [DEBIT:0] score_8_x30;
wire signed [DEBIT:0] score_8_x31;
wire signed [DEBIT:0] score_8_x32;
wire signed [DEBIT:0] score_8_x33;
wire signed [DEBIT:0] score_8_x34;
wire signed [DEBIT:0] score_8_x35;
wire signed [DEBIT:0] score_8_x36;
wire signed [DEBIT:0] score_8_x37;
wire signed [DEBIT:0] score_8_x38;
wire signed [DEBIT:0] score_8_x39;
wire signed [DEBIT:0] score_8_x40;
wire signed [DEBIT:0] score_8_x41;
wire signed [DEBIT:0] score_8_x42;
wire signed [DEBIT:0] score_8_x43;
wire signed [DEBIT:0] score_8_x44;
wire signed [DEBIT:0] score_8_x45;
wire signed [DEBIT:0] score_8_x46;
wire signed [DEBIT:0] score_8_x47;
wire signed [DEBIT:0] score_8_x48;
wire signed [DEBIT:0] score_8_x49;
wire signed [DEBIT:0] score_8_x50;
wire signed [DEBIT:0] score_8_x51;
wire signed [DEBIT:0] score_8_x52;
wire signed [DEBIT:0] score_8_x53;
wire signed [DEBIT:0] score_8_x54;
wire signed [DEBIT:0] score_8_x55;
wire signed [DEBIT:0] score_8_x56;
wire signed [DEBIT:0] score_8_x57;
wire signed [DEBIT:0] score_8_x58;
wire signed [DEBIT:0] score_8_x59;
wire signed [DEBIT:0] score_8_x60;
wire signed [DEBIT:0] score_8_x61;
wire signed [DEBIT:0] score_8_x62;
wire signed [DEBIT:0] score_8_x63;
wire signed [DEBIT:0] score_8_x64;
wire signed [DEBIT:0] score_8_x65;
wire signed [DEBIT:0] score_8_x66;
wire signed [DEBIT:0] score_8_x67;
wire signed [DEBIT:0] score_8_x68;
wire signed [DEBIT:0] score_8_x69;
wire signed [DEBIT:0] score_8_x70;
wire signed [DEBIT:0] score_8_x71;
wire signed [DEBIT:0] score_8_x72;
wire signed [DEBIT:0] score_8_x73;
wire signed [DEBIT:0] score_8_x74;
wire signed [DEBIT:0] score_8_x75;
wire signed [DEBIT:0] score_8_x76;
wire signed [DEBIT:0] score_8_x77;
wire signed [DEBIT:0] score_8_x78;
wire signed [DEBIT:0] score_8_x79;
wire signed [DEBIT:0] score_8_x80;
wire signed [DEBIT:0] score_8_x81;
wire signed [DEBIT:0] score_8_x82;
wire signed [DEBIT:0] score_8_x83;
wire signed [DEBIT:0] score_8_x84;
wire signed [DEBIT:0] score_8_x85;
wire signed [DEBIT:0] score_8_x86;
wire signed [DEBIT:0] score_8_x87;
wire signed [DEBIT:0] score_8_x88;
wire signed [DEBIT:0] score_8_x89;
wire signed [DEBIT:0] score_8_x90;
wire signed [DEBIT:0] score_8_x91;
wire signed [DEBIT:0] score_8_x92;
wire signed [DEBIT:0] score_8_x93;
wire signed [DEBIT:0] score_8_x94;
wire signed [DEBIT:0] score_8_x95;
wire signed [DEBIT:0] score_8_x96;
wire signed [DEBIT:0] score_8_x97;
wire signed [DEBIT:0] score_8_x98;
wire signed [DEBIT:0] score_8_x99;
wire signed [DEBIT:0] score_8_x100;
wire signed [DEBIT:0] score_8_x101;
wire signed [DEBIT:0] score_8_x102;
wire signed [DEBIT:0] score_8_x103;
wire signed [DEBIT:0] score_8_x104;
wire signed [DEBIT:0] score_8_x105;
wire signed [DEBIT:0] score_8_x106;
wire signed [DEBIT:0] score_8_x107;
wire signed [DEBIT:0] score_8_x108;
wire signed [DEBIT:0] score_8_x109;
wire signed [DEBIT:0] score_8_x110;
wire signed [DEBIT:0] score_8_x111;
wire signed [DEBIT:0] score_8_x112;
wire signed [DEBIT:0] score_8_x113;
wire signed [DEBIT:0] score_8_x114;
wire signed [DEBIT:0] score_8_x115;
wire signed [DEBIT:0] score_8_x116;
wire signed [DEBIT:0] score_8_x117;
wire signed [DEBIT:0] score_8_x118;
wire signed [DEBIT:0] score_8_x119;
wire signed [DEBIT:0] score_8_x120;
wire signed [DEBIT:0] score_8_x121;
wire signed [DEBIT:0] score_8_x122;
wire signed [DEBIT:0] score_8_x123;
wire signed [DEBIT:0] score_8_x124;
wire signed [DEBIT:0] score_8_x125;
wire signed [DEBIT:0] score_8_x126;
wire signed [DEBIT:0] score_8_x127;
wire signed [DEBIT:0] score_8_x128;
wire signed [DEBIT:0] score_8_x129;
wire signed [DEBIT:0] score_8_x130;
wire signed [DEBIT:0] score_8_x131;
wire signed [DEBIT:0] score_8_x132;
wire signed [DEBIT:0] score_8_x133;
wire signed [DEBIT:0] score_8_x134;
wire signed [DEBIT:0] score_8_x135;
wire signed [DEBIT:0] score_8_x136;
wire signed [DEBIT:0] score_8_x137;
wire signed [DEBIT:0] score_8_x138;
wire signed [DEBIT:0] score_8_x139;
wire signed [DEBIT:0] score_8_x140;
wire signed [DEBIT:0] score_8_x141;
wire signed [DEBIT:0] score_8_x142;
wire signed [DEBIT:0] score_8_x143;
wire signed [DEBIT:0] score_8_x144;
wire signed [DEBIT:0] score_8_x145;
wire signed [DEBIT:0] score_8_x146;
wire signed [DEBIT:0] score_8_x147;
wire signed [DEBIT:0] score_8_x148;
wire signed [DEBIT:0] score_8_x149;
wire signed [DEBIT:0] score_8_x150;
wire signed [DEBIT:0] score_8_x151;
wire signed [DEBIT:0] score_8_x152;
wire signed [DEBIT:0] score_8_x153;
wire signed [DEBIT:0] score_8_x154;
wire signed [DEBIT:0] score_8_x155;
wire signed [DEBIT:0] score_8_x156;
wire signed [DEBIT:0] score_8_x157;
wire signed [DEBIT:0] score_8_x158;
wire signed [DEBIT:0] score_8_x159;
wire signed [DEBIT:0] score_8_x160;
wire signed [DEBIT:0] score_8_x161;
wire signed [DEBIT:0] score_8_x162;
wire signed [DEBIT:0] score_8_x163;
wire signed [DEBIT:0] score_8_x164;
wire signed [DEBIT:0] score_8_x165;
wire signed [DEBIT:0] score_8_x166;
wire signed [DEBIT:0] score_8_x167;
wire signed [DEBIT:0] score_8_x168;
wire signed [DEBIT:0] score_8_x169;
wire signed [DEBIT:0] score_8_x170;
wire signed [DEBIT:0] score_8_x171;
wire signed [DEBIT:0] score_8_x172;
wire signed [DEBIT:0] score_8_x173;
wire signed [DEBIT:0] score_8_x174;
wire signed [DEBIT:0] score_8_x175;
wire signed [DEBIT:0] score_8_x176;
wire signed [DEBIT:0] score_8_x177;
wire signed [DEBIT:0] score_8_x178;
wire signed [DEBIT:0] score_8_x179;
wire signed [DEBIT:0] score_8_x180;
wire signed [DEBIT:0] score_8_x181;
wire signed [DEBIT:0] score_8_x182;
wire signed [DEBIT:0] score_8_x183;
wire signed [DEBIT:0] score_8_x184;
wire signed [DEBIT:0] score_8_x185;
wire signed [DEBIT:0] score_8_x186;
wire signed [DEBIT:0] score_8_x187;
wire signed [DEBIT:0] score_8_x188;
wire signed [DEBIT:0] score_8_x189;
wire signed [DEBIT:0] score_8_x190;
wire signed [DEBIT:0] score_8_x191;
wire signed [DEBIT:0] score_8_x192;
wire signed [DEBIT:0] score_8_x193;
wire signed [DEBIT:0] score_8_x194;
wire signed [DEBIT:0] score_8_x195;
wire signed [DEBIT:0] score_8_x196;
wire signed [DEBIT:0] score_8_x197;
wire signed [DEBIT:0] score_8_x198;
wire signed [DEBIT:0] score_8_x199;
wire signed [DEBIT:0] score_8_x200;
wire signed [DEBIT:0] score_8_x201;
wire signed [DEBIT:0] score_8_x202;
wire signed [DEBIT:0] score_8_x203;
wire signed [DEBIT:0] score_8_x204;
wire signed [DEBIT:0] score_8_x205;
wire signed [DEBIT:0] score_8_x206;
wire signed [DEBIT:0] score_8_x207;
wire signed [DEBIT:0] score_8_x208;
wire signed [DEBIT:0] score_8_x209;
wire signed [DEBIT:0] score_8_x210;
wire signed [DEBIT:0] score_8_x211;
wire signed [DEBIT:0] score_8_x212;
wire signed [DEBIT:0] score_8_x213;
wire signed [DEBIT:0] score_8_x214;
wire signed [DEBIT:0] score_8_x215;
wire signed [DEBIT:0] score_8_x216;
wire signed [DEBIT:0] score_8_x217;
wire signed [DEBIT:0] score_8_x218;
wire signed [DEBIT:0] score_8_x219;
wire signed [DEBIT:0] score_8_x220;
wire signed [DEBIT:0] score_8_x221;
wire signed [DEBIT:0] score_8_x222;
wire signed [DEBIT:0] score_8_x223;
wire signed [DEBIT:0] score_8_x224;
wire signed [DEBIT:0] score_8_x225;
wire signed [DEBIT:0] score_8_x226;
wire signed [DEBIT:0] score_8_x227;
wire signed [DEBIT:0] score_8_x228;
wire signed [DEBIT:0] score_8_x229;
wire signed [DEBIT:0] score_8_x230;
wire signed [DEBIT:0] score_8_x231;
wire signed [DEBIT:0] score_8_x232;
wire signed [DEBIT:0] score_8_x233;
wire signed [DEBIT:0] score_8_x234;
wire signed [DEBIT:0] score_8_x235;
wire signed [DEBIT:0] score_8_x236;
wire signed [DEBIT:0] score_8_x237;
wire signed [DEBIT:0] score_8_x238;
wire signed [DEBIT:0] score_8_x239;
wire signed [DEBIT:0] score_8_x240;
wire signed [DEBIT:0] score_8_x241;
wire signed [DEBIT:0] score_8_x242;
wire signed [DEBIT:0] score_8_x243;
wire signed [DEBIT:0] score_8_x244;
wire signed [DEBIT:0] score_8_x245;
wire signed [DEBIT:0] score_8_x246;
wire signed [DEBIT:0] score_8_x247;
wire signed [DEBIT:0] score_8_x248;
wire signed [DEBIT:0] score_8_x249;
wire signed [DEBIT:0] score_8_x250;
wire signed [DEBIT:0] score_8_x251;
wire signed [DEBIT:0] score_8_x252;
wire signed [DEBIT:0] score_8_x253;
wire signed [DEBIT:0] score_8_x254;
wire signed [DEBIT:0] score_8_x255;
wire signed [DEBIT:0] score_8_x256;
wire signed [DEBIT:0] score_8_x257;
wire signed [DEBIT:0] score_8_x258;
wire signed [DEBIT:0] score_8_x259;
wire signed [DEBIT:0] score_8_x260;
wire signed [DEBIT:0] score_8_x261;
wire signed [DEBIT:0] score_8_x262;
wire signed [DEBIT:0] score_8_x263;
wire signed [DEBIT:0] score_8_x264;
wire signed [DEBIT:0] score_8_x265;
wire signed [DEBIT:0] score_8_x266;
wire signed [DEBIT:0] score_8_x267;
wire signed [DEBIT:0] score_8_x268;
wire signed [DEBIT:0] score_8_x269;
wire signed [DEBIT:0] score_8_x270;
wire signed [DEBIT:0] score_8_x271;
wire signed [DEBIT:0] score_8_x272;
wire signed [DEBIT:0] score_8_x273;
wire signed [DEBIT:0] score_8_x274;
wire signed [DEBIT:0] score_8_x275;
wire signed [DEBIT:0] score_8_x276;
wire signed [DEBIT:0] score_8_x277;
wire signed [DEBIT:0] score_8_x278;
wire signed [DEBIT:0] score_8_x279;
wire signed [DEBIT:0] score_8_x280;
wire signed [DEBIT:0] score_8_x281;
wire signed [DEBIT:0] score_8_x282;
wire signed [DEBIT:0] score_8_x283;
wire signed [DEBIT:0] score_8_x284;
wire signed [DEBIT:0] score_8_x285;
wire signed [DEBIT:0] score_8_x286;
wire signed [DEBIT:0] score_8_x287;
wire signed [DEBIT:0] score_8_x288;
wire signed [DEBIT:0] score_8_x289;
wire signed [DEBIT:0] score_8_x290;
wire signed [DEBIT:0] score_8_x291;
wire signed [DEBIT:0] score_8_x292;
wire signed [DEBIT:0] score_8_x293;
wire signed [DEBIT:0] score_8_x294;
wire signed [DEBIT:0] score_8_x295;
wire signed [DEBIT:0] score_8_x296;
wire signed [DEBIT:0] score_8_x297;
wire signed [DEBIT:0] score_8_x298;
wire signed [DEBIT:0] score_8_x299;
wire signed [DEBIT:0] score_8_x300;
wire signed [DEBIT:0] score_8_x301;
wire signed [DEBIT:0] score_8_x302;
wire signed [DEBIT:0] score_8_x303;
wire signed [DEBIT:0] score_8_x304;
wire signed [DEBIT:0] score_8_x305;
wire signed [DEBIT:0] score_8_x306;
wire signed [DEBIT:0] score_8_x307;
wire signed [DEBIT:0] score_8_x308;
wire signed [DEBIT:0] score_8_x309;
wire signed [DEBIT:0] score_8_x310;
wire signed [DEBIT:0] score_8_x311;
wire signed [DEBIT:0] score_8_x312;
wire signed [DEBIT:0] score_8_x313;
wire signed [DEBIT:0] score_8_x314;
wire signed [DEBIT:0] score_8_x315;
wire signed [DEBIT:0] score_8_x316;
wire signed [DEBIT:0] score_8_x317;
wire signed [DEBIT:0] score_8_x318;
wire signed [DEBIT:0] score_8_x319;
wire signed [DEBIT:0] score_8_x320;
wire signed [DEBIT:0] score_8_x321;
wire signed [DEBIT:0] score_8_x322;
wire signed [DEBIT:0] score_8_x323;
wire signed [DEBIT:0] score_8_x324;
wire signed [DEBIT:0] score_8_x325;
wire signed [DEBIT:0] score_8_x326;
wire signed [DEBIT:0] score_8_x327;
wire signed [DEBIT:0] score_8_x328;
wire signed [DEBIT:0] score_8_x329;
wire signed [DEBIT:0] score_8_x330;
wire signed [DEBIT:0] score_8_x331;
wire signed [DEBIT:0] score_8_x332;
wire signed [DEBIT:0] score_8_x333;
wire signed [DEBIT:0] score_8_x334;
wire signed [DEBIT:0] score_8_x335;
wire signed [DEBIT:0] score_8_x336;
wire signed [DEBIT:0] score_8_x337;
wire signed [DEBIT:0] score_8_x338;
wire signed [DEBIT:0] score_8_x339;
wire signed [DEBIT:0] score_8_x340;
wire signed [DEBIT:0] score_8_x341;
wire signed [DEBIT:0] score_8_x342;
wire signed [DEBIT:0] score_8_x343;
wire signed [DEBIT:0] score_8_x344;
wire signed [DEBIT:0] score_8_x345;
wire signed [DEBIT:0] score_8_x346;
wire signed [DEBIT:0] score_8_x347;
wire signed [DEBIT:0] score_8_x348;
wire signed [DEBIT:0] score_8_x349;
wire signed [DEBIT:0] score_8_x350;
wire signed [DEBIT:0] score_8_x351;
wire signed [DEBIT:0] score_8_x352;
wire signed [DEBIT:0] score_8_x353;
wire signed [DEBIT:0] score_8_x354;
wire signed [DEBIT:0] score_8_x355;
wire signed [DEBIT:0] score_8_x356;
wire signed [DEBIT:0] score_8_x357;
wire signed [DEBIT:0] score_8_x358;
wire signed [DEBIT:0] score_8_x359;
wire signed [DEBIT:0] score_8_x360;
wire signed [DEBIT:0] score_8_x361;
wire signed [DEBIT:0] score_8_x362;
wire signed [DEBIT:0] score_8_x363;
wire signed [DEBIT:0] score_8_x364;
wire signed [DEBIT:0] score_8_x365;
wire signed [DEBIT:0] score_8_x366;
wire signed [DEBIT:0] score_8_x367;
wire signed [DEBIT:0] score_8_x368;
wire signed [DEBIT:0] score_8_x369;
wire signed [DEBIT:0] score_8_x370;
wire signed [DEBIT:0] score_8_x371;
wire signed [DEBIT:0] score_8_x372;
wire signed [DEBIT:0] score_8_x373;
wire signed [DEBIT:0] score_8_x374;
wire signed [DEBIT:0] score_8_x375;
wire signed [DEBIT:0] score_8_x376;
wire signed [DEBIT:0] score_8_x377;
wire signed [DEBIT:0] score_8_x378;
wire signed [DEBIT:0] score_8_x379;
wire signed [DEBIT:0] score_8_x380;
wire signed [DEBIT:0] score_8_x381;
wire signed [DEBIT:0] score_8_x382;
wire signed [DEBIT:0] score_8_x383;
wire signed [DEBIT:0] score_8_x384;
wire signed [DEBIT:0] score_8_x385;
wire signed [DEBIT:0] score_8_x386;
wire signed [DEBIT:0] score_8_x387;
wire signed [DEBIT:0] score_8_x388;
wire signed [DEBIT:0] score_8_x389;
wire signed [DEBIT:0] score_8_x390;
wire signed [DEBIT:0] score_8_x391;
wire signed [DEBIT:0] score_8_x392;
wire signed [DEBIT:0] score_8_x393;
wire signed [DEBIT:0] score_8_x394;
wire signed [DEBIT:0] score_8_x395;
wire signed [DEBIT:0] score_8_x396;
wire signed [DEBIT:0] score_8_x397;
wire signed [DEBIT:0] score_8_x398;
wire signed [DEBIT:0] score_8_x399;
wire signed [DEBIT:0] score_8_x400;
wire signed [DEBIT:0] score_8_x401;
wire signed [DEBIT:0] score_8_x402;
wire signed [DEBIT:0] score_8_x403;
wire signed [DEBIT:0] score_8_x404;
wire signed [DEBIT:0] score_8_x405;
wire signed [DEBIT:0] score_8_x406;
wire signed [DEBIT:0] score_8_x407;
wire signed [DEBIT:0] score_8_x408;
wire signed [DEBIT:0] score_8_x409;
wire signed [DEBIT:0] score_8_x410;
wire signed [DEBIT:0] score_8_x411;
wire signed [DEBIT:0] score_8_x412;
wire signed [DEBIT:0] score_8_x413;
wire signed [DEBIT:0] score_8_x414;
wire signed [DEBIT:0] score_8_x415;
wire signed [DEBIT:0] score_8_x416;
wire signed [DEBIT:0] score_8_x417;
wire signed [DEBIT:0] score_8_x418;
wire signed [DEBIT:0] score_8_x419;
wire signed [DEBIT:0] score_8_x420;
wire signed [DEBIT:0] score_8_x421;
wire signed [DEBIT:0] score_8_x422;
wire signed [DEBIT:0] score_8_x423;
wire signed [DEBIT:0] score_8_x424;
wire signed [DEBIT:0] score_8_x425;
wire signed [DEBIT:0] score_8_x426;
wire signed [DEBIT:0] score_8_x427;
wire signed [DEBIT:0] score_8_x428;
wire signed [DEBIT:0] score_8_x429;
wire signed [DEBIT:0] score_8_x430;
wire signed [DEBIT:0] score_8_x431;
wire signed [DEBIT:0] score_8_x432;
wire signed [DEBIT:0] score_8_x433;
wire signed [DEBIT:0] score_8_x434;
wire signed [DEBIT:0] score_8_x435;
wire signed [DEBIT:0] score_8_x436;
wire signed [DEBIT:0] score_8_x437;
wire signed [DEBIT:0] score_8_x438;
wire signed [DEBIT:0] score_8_x439;
wire signed [DEBIT:0] score_8_x440;
wire signed [DEBIT:0] score_8_x441;
wire signed [DEBIT:0] score_8_x442;
wire signed [DEBIT:0] score_8_x443;
wire signed [DEBIT:0] score_8_x444;
wire signed [DEBIT:0] score_8_x445;
wire signed [DEBIT:0] score_8_x446;
wire signed [DEBIT:0] score_8_x447;
wire signed [DEBIT:0] score_8_x448;
wire signed [DEBIT:0] score_8_x449;
wire signed [DEBIT:0] score_8_x450;
wire signed [DEBIT:0] score_8_x451;
wire signed [DEBIT:0] score_8_x452;
wire signed [DEBIT:0] score_8_x453;
wire signed [DEBIT:0] score_8_x454;
wire signed [DEBIT:0] score_8_x455;
wire signed [DEBIT:0] score_8_x456;
wire signed [DEBIT:0] score_8_x457;
wire signed [DEBIT:0] score_8_x458;
wire signed [DEBIT:0] score_8_x459;
wire signed [DEBIT:0] score_8_x460;
wire signed [DEBIT:0] score_8_x461;
wire signed [DEBIT:0] score_8_x462;
wire signed [DEBIT:0] score_8_x463;
wire signed [DEBIT:0] score_8_x464;
wire signed [DEBIT:0] score_8_x465;
wire signed [DEBIT:0] score_8_x466;
wire signed [DEBIT:0] score_8_x467;
wire signed [DEBIT:0] score_8_x468;
wire signed [DEBIT:0] score_8_x469;
wire signed [DEBIT:0] score_8_x470;
wire signed [DEBIT:0] score_8_x471;
wire signed [DEBIT:0] score_8_x472;
wire signed [DEBIT:0] score_8_x473;
wire signed [DEBIT:0] score_8_x474;
wire signed [DEBIT:0] score_8_x475;
wire signed [DEBIT:0] score_8_x476;
wire signed [DEBIT:0] score_8_x477;
wire signed [DEBIT:0] score_8_x478;
wire signed [DEBIT:0] score_8_x479;
wire signed [DEBIT:0] score_8_x480;
wire signed [DEBIT:0] score_8_x481;
wire signed [DEBIT:0] score_8_x482;
wire signed [DEBIT:0] score_8_x483;
wire signed [DEBIT:0] score_8_x484;
wire signed [DEBIT:0] score_8_x485;
wire signed [DEBIT:0] score_8_x486;
wire signed [DEBIT:0] score_8_x487;
wire signed [DEBIT:0] score_8_x488;
wire signed [DEBIT:0] score_8_x489;
wire signed [DEBIT:0] score_8_x490;
wire signed [DEBIT:0] score_8_x491;
wire signed [DEBIT:0] score_8_x492;
wire signed [DEBIT:0] score_8_x493;
wire signed [DEBIT:0] score_8_x494;
wire signed [DEBIT:0] score_8_x495;
wire signed [DEBIT:0] score_8_x496;
wire signed [DEBIT:0] score_8_x497;
wire signed [DEBIT:0] score_8_x498;
wire signed [DEBIT:0] score_8_x499;
wire signed [DEBIT:0] score_8_x500;
wire signed [DEBIT:0] score_8_x501;
wire signed [DEBIT:0] score_8_x502;
wire signed [DEBIT:0] score_8_x503;
wire signed [DEBIT:0] score_8_x504;
wire signed [DEBIT:0] score_8_x505;
wire signed [DEBIT:0] score_8_x506;
wire signed [DEBIT:0] score_8_x507;
wire signed [DEBIT:0] score_8_x508;
wire signed [DEBIT:0] score_8_x509;
wire signed [DEBIT:0] score_8_x510;
wire signed [DEBIT:0] score_8_x511;
wire signed [DEBIT:0] score_8_x512;
wire signed [DEBIT:0] score_8_x513;
wire signed [DEBIT:0] score_8_x514;
wire signed [DEBIT:0] score_8_x515;
wire signed [DEBIT:0] score_8_x516;
wire signed [DEBIT:0] score_8_x517;
wire signed [DEBIT:0] score_8_x518;
wire signed [DEBIT:0] score_8_x519;
wire signed [DEBIT:0] score_8_x520;
wire signed [DEBIT:0] score_8_x521;
wire signed [DEBIT:0] score_8_x522;
wire signed [DEBIT:0] score_8_x523;
wire signed [DEBIT:0] score_8_x524;
wire signed [DEBIT:0] score_8_x525;
wire signed [DEBIT:0] score_8_x526;
wire signed [DEBIT:0] score_8_x527;
wire signed [DEBIT:0] score_8_x528;
wire signed [DEBIT:0] score_8_x529;
wire signed [DEBIT:0] score_8_x530;
wire signed [DEBIT:0] score_8_x531;
wire signed [DEBIT:0] score_8_x532;
wire signed [DEBIT:0] score_8_x533;
wire signed [DEBIT:0] score_8_x534;
wire signed [DEBIT:0] score_8_x535;
wire signed [DEBIT:0] score_8_x536;
wire signed [DEBIT:0] score_8_x537;
wire signed [DEBIT:0] score_8_x538;
wire signed [DEBIT:0] score_8_x539;
wire signed [DEBIT:0] score_8_x540;
wire signed [DEBIT:0] score_8_x541;
wire signed [DEBIT:0] score_8_x542;
wire signed [DEBIT:0] score_8_x543;
wire signed [DEBIT:0] score_8_x544;
wire signed [DEBIT:0] score_8_x545;
wire signed [DEBIT:0] score_8_x546;
wire signed [DEBIT:0] score_8_x547;
wire signed [DEBIT:0] score_8_x548;
wire signed [DEBIT:0] score_8_x549;
wire signed [DEBIT:0] score_8_x550;
wire signed [DEBIT:0] score_8_x551;
wire signed [DEBIT:0] score_8_x552;
wire signed [DEBIT:0] score_8_x553;
wire signed [DEBIT:0] score_8_x554;
wire signed [DEBIT:0] score_8_x555;
wire signed [DEBIT:0] score_8_x556;
wire signed [DEBIT:0] score_8_x557;
wire signed [DEBIT:0] score_8_x558;
wire signed [DEBIT:0] score_8_x559;
wire signed [DEBIT:0] score_8_x560;
wire signed [DEBIT:0] score_8_x561;
wire signed [DEBIT:0] score_8_x562;
wire signed [DEBIT:0] score_8_x563;
wire signed [DEBIT:0] score_8_x564;
wire signed [DEBIT:0] score_8_x565;
wire signed [DEBIT:0] score_8_x566;
wire signed [DEBIT:0] score_8_x567;
wire signed [DEBIT:0] score_8_x568;
wire signed [DEBIT:0] score_8_x569;
wire signed [DEBIT:0] score_8_x570;
wire signed [DEBIT:0] score_8_x571;
wire signed [DEBIT:0] score_8_x572;
wire signed [DEBIT:0] score_8_x573;
wire signed [DEBIT:0] score_8_x574;
wire signed [DEBIT:0] score_8_x575;
wire signed [DEBIT:0] score_8_x576;
wire signed [DEBIT:0] score_8_x577;
wire signed [DEBIT:0] score_8_x578;
wire signed [DEBIT:0] score_8_x579;
wire signed [DEBIT:0] score_8_x580;
wire signed [DEBIT:0] score_8_x581;
wire signed [DEBIT:0] score_8_x582;
wire signed [DEBIT:0] score_8_x583;
wire signed [DEBIT:0] score_8_x584;
wire signed [DEBIT:0] score_8_x585;
wire signed [DEBIT:0] score_8_x586;
wire signed [DEBIT:0] score_8_x587;
wire signed [DEBIT:0] score_8_x588;
wire signed [DEBIT:0] score_8_x589;
wire signed [DEBIT:0] score_8_x590;
wire signed [DEBIT:0] score_8_x591;
wire signed [DEBIT:0] score_8_x592;
wire signed [DEBIT:0] score_8_x593;
wire signed [DEBIT:0] score_8_x594;
wire signed [DEBIT:0] score_8_x595;
wire signed [DEBIT:0] score_8_x596;
wire signed [DEBIT:0] score_8_x597;
wire signed [DEBIT:0] score_8_x598;
wire signed [DEBIT:0] score_8_x599;
wire signed [DEBIT:0] score_8_x600;
wire signed [DEBIT:0] score_8_x601;
wire signed [DEBIT:0] score_8_x602;
wire signed [DEBIT:0] score_8_x603;
wire signed [DEBIT:0] score_8_x604;
wire signed [DEBIT:0] score_8_x605;
wire signed [DEBIT:0] score_8_x606;
wire signed [DEBIT:0] score_8_x607;
wire signed [DEBIT:0] score_8_x608;
wire signed [DEBIT:0] score_8_x609;
wire signed [DEBIT:0] score_8_x610;
wire signed [DEBIT:0] score_8_x611;
wire signed [DEBIT:0] score_8_x612;
wire signed [DEBIT:0] score_8_x613;
wire signed [DEBIT:0] score_8_x614;
wire signed [DEBIT:0] score_8_x615;
wire signed [DEBIT:0] score_8_x616;
wire signed [DEBIT:0] score_8_x617;
wire signed [DEBIT:0] score_8_x618;
wire signed [DEBIT:0] score_8_x619;
wire signed [DEBIT:0] score_8_x620;
wire signed [DEBIT:0] score_8_x621;
wire signed [DEBIT:0] score_8_x622;
wire signed [DEBIT:0] score_8_x623;
wire signed [DEBIT:0] score_8_x624;
wire signed [DEBIT:0] score_8_x625;
wire signed [DEBIT:0] score_8_x626;
wire signed [DEBIT:0] score_8_x627;
wire signed [DEBIT:0] score_8_x628;
wire signed [DEBIT:0] score_8_x629;
wire signed [DEBIT:0] score_8_x630;
wire signed [DEBIT:0] score_8_x631;
wire signed [DEBIT:0] score_8_x632;
wire signed [DEBIT:0] score_8_x633;
wire signed [DEBIT:0] score_8_x634;
wire signed [DEBIT:0] score_8_x635;
wire signed [DEBIT:0] score_8_x636;
wire signed [DEBIT:0] score_8_x637;
wire signed [DEBIT:0] score_8_x638;
wire signed [DEBIT:0] score_8_x639;
wire signed [DEBIT:0] score_8_x640;
wire signed [DEBIT:0] score_8_x641;
wire signed [DEBIT:0] score_8_x642;
wire signed [DEBIT:0] score_8_x643;
wire signed [DEBIT:0] score_8_x644;
wire signed [DEBIT:0] score_8_x645;
wire signed [DEBIT:0] score_8_x646;
wire signed [DEBIT:0] score_8_x647;
wire signed [DEBIT:0] score_8_x648;
wire signed [DEBIT:0] score_8_x649;
wire signed [DEBIT:0] score_8_x650;
wire signed [DEBIT:0] score_8_x651;
wire signed [DEBIT:0] score_8_x652;
wire signed [DEBIT:0] score_8_x653;
wire signed [DEBIT:0] score_8_x654;
wire signed [DEBIT:0] score_8_x655;
wire signed [DEBIT:0] score_8_x656;
wire signed [DEBIT:0] score_8_x657;
wire signed [DEBIT:0] score_8_x658;
wire signed [DEBIT:0] score_8_x659;
wire signed [DEBIT:0] score_8_x660;
wire signed [DEBIT:0] score_8_x661;
wire signed [DEBIT:0] score_8_x662;
wire signed [DEBIT:0] score_8_x663;
wire signed [DEBIT:0] score_8_x664;
wire signed [DEBIT:0] score_8_x665;
wire signed [DEBIT:0] score_8_x666;
wire signed [DEBIT:0] score_8_x667;
wire signed [DEBIT:0] score_8_x668;
wire signed [DEBIT:0] score_8_x669;
wire signed [DEBIT:0] score_8_x670;
wire signed [DEBIT:0] score_8_x671;
wire signed [DEBIT:0] score_8_x672;
wire signed [DEBIT:0] score_8_x673;
wire signed [DEBIT:0] score_8_x674;
wire signed [DEBIT:0] score_8_x675;
wire signed [DEBIT:0] score_8_x676;
wire signed [DEBIT:0] score_8_x677;
wire signed [DEBIT:0] score_8_x678;
wire signed [DEBIT:0] score_8_x679;
wire signed [DEBIT:0] score_8_x680;
wire signed [DEBIT:0] score_8_x681;
wire signed [DEBIT:0] score_8_x682;
wire signed [DEBIT:0] score_8_x683;
wire signed [DEBIT:0] score_8_x684;
wire signed [DEBIT:0] score_8_x685;
wire signed [DEBIT:0] score_8_x686;
wire signed [DEBIT:0] score_8_x687;
wire signed [DEBIT:0] score_8_x688;
wire signed [DEBIT:0] score_8_x689;
wire signed [DEBIT:0] score_8_x690;
wire signed [DEBIT:0] score_8_x691;
wire signed [DEBIT:0] score_8_x692;
wire signed [DEBIT:0] score_8_x693;
wire signed [DEBIT:0] score_8_x694;
wire signed [DEBIT:0] score_8_x695;
wire signed [DEBIT:0] score_8_x696;
wire signed [DEBIT:0] score_8_x697;
wire signed [DEBIT:0] score_8_x698;
wire signed [DEBIT:0] score_8_x699;
wire signed [DEBIT:0] score_8_x700;
wire signed [DEBIT:0] score_8_x701;
wire signed [DEBIT:0] score_8_x702;
wire signed [DEBIT:0] score_8_x703;
wire signed [DEBIT:0] score_8_x704;
wire signed [DEBIT:0] score_8_x705;
wire signed [DEBIT:0] score_8_x706;
wire signed [DEBIT:0] score_8_x707;
wire signed [DEBIT:0] score_8_x708;
wire signed [DEBIT:0] score_8_x709;
wire signed [DEBIT:0] score_8_x710;
wire signed [DEBIT:0] score_8_x711;
wire signed [DEBIT:0] score_8_x712;
wire signed [DEBIT:0] score_8_x713;
wire signed [DEBIT:0] score_8_x714;
wire signed [DEBIT:0] score_8_x715;
wire signed [DEBIT:0] score_8_x716;
wire signed [DEBIT:0] score_8_x717;
wire signed [DEBIT:0] score_8_x718;
wire signed [DEBIT:0] score_8_x719;
wire signed [DEBIT:0] score_8_x720;
wire signed [DEBIT:0] score_8_x721;
wire signed [DEBIT:0] score_8_x722;
wire signed [DEBIT:0] score_8_x723;
wire signed [DEBIT:0] score_8_x724;
wire signed [DEBIT:0] score_8_x725;
wire signed [DEBIT:0] score_8_x726;
wire signed [DEBIT:0] score_8_x727;
wire signed [DEBIT:0] score_8_x728;
wire signed [DEBIT:0] score_8_x729;
wire signed [DEBIT:0] score_8_x730;
wire signed [DEBIT:0] score_8_x731;
wire signed [DEBIT:0] score_8_x732;
wire signed [DEBIT:0] score_8_x733;
wire signed [DEBIT:0] score_8_x734;
wire signed [DEBIT:0] score_8_x735;
wire signed [DEBIT:0] score_8_x736;
wire signed [DEBIT:0] score_8_x737;
wire signed [DEBIT:0] score_8_x738;
wire signed [DEBIT:0] score_8_x739;
wire signed [DEBIT:0] score_8_x740;
wire signed [DEBIT:0] score_8_x741;
wire signed [DEBIT:0] score_8_x742;
wire signed [DEBIT:0] score_8_x743;
wire signed [DEBIT:0] score_8_x744;
wire signed [DEBIT:0] score_8_x745;
wire signed [DEBIT:0] score_8_x746;
wire signed [DEBIT:0] score_8_x747;
wire signed [DEBIT:0] score_8_x748;
wire signed [DEBIT:0] score_8_x749;
wire signed [DEBIT:0] score_8_x750;
wire signed [DEBIT:0] score_8_x751;
wire signed [DEBIT:0] score_8_x752;
wire signed [DEBIT:0] score_8_x753;
wire signed [DEBIT:0] score_8_x754;
wire signed [DEBIT:0] score_8_x755;
wire signed [DEBIT:0] score_8_x756;
wire signed [DEBIT:0] score_8_x757;
wire signed [DEBIT:0] score_8_x758;
wire signed [DEBIT:0] score_8_x759;
wire signed [DEBIT:0] score_8_x760;
wire signed [DEBIT:0] score_8_x761;
wire signed [DEBIT:0] score_8_x762;
wire signed [DEBIT:0] score_8_x763;
wire signed [DEBIT:0] score_8_x764;
wire signed [DEBIT:0] score_8_x765;
wire signed [DEBIT:0] score_8_x766;
wire signed [DEBIT:0] score_8_x767;
wire signed [DEBIT:0] score_8_x768;
wire signed [DEBIT:0] score_8_x769;
wire signed [DEBIT:0] score_8_x770;
wire signed [DEBIT:0] score_8_x771;
wire signed [DEBIT:0] score_8_x772;
wire signed [DEBIT:0] score_8_x773;
wire signed [DEBIT:0] score_8_x774;
wire signed [DEBIT:0] score_8_x775;
wire signed [DEBIT:0] score_8_x776;
wire signed [DEBIT:0] score_8_x777;
wire signed [DEBIT:0] score_8_x778;
wire signed [DEBIT:0] score_8_x779;
wire signed [DEBIT:0] score_8_x780;
wire signed [DEBIT:0] score_8_x781;
wire signed [DEBIT:0] score_8_x782;
wire signed [DEBIT:0] score_8_x783;
wire signed [DEBIT:0] score_8_x784;
wire signed [DEBIT:0] score_9_x1;
wire signed [DEBIT:0] score_9_x2;
wire signed [DEBIT:0] score_9_x3;
wire signed [DEBIT:0] score_9_x4;
wire signed [DEBIT:0] score_9_x5;
wire signed [DEBIT:0] score_9_x6;
wire signed [DEBIT:0] score_9_x7;
wire signed [DEBIT:0] score_9_x8;
wire signed [DEBIT:0] score_9_x9;
wire signed [DEBIT:0] score_9_x10;
wire signed [DEBIT:0] score_9_x11;
wire signed [DEBIT:0] score_9_x12;
wire signed [DEBIT:0] score_9_x13;
wire signed [DEBIT:0] score_9_x14;
wire signed [DEBIT:0] score_9_x15;
wire signed [DEBIT:0] score_9_x16;
wire signed [DEBIT:0] score_9_x17;
wire signed [DEBIT:0] score_9_x18;
wire signed [DEBIT:0] score_9_x19;
wire signed [DEBIT:0] score_9_x20;
wire signed [DEBIT:0] score_9_x21;
wire signed [DEBIT:0] score_9_x22;
wire signed [DEBIT:0] score_9_x23;
wire signed [DEBIT:0] score_9_x24;
wire signed [DEBIT:0] score_9_x25;
wire signed [DEBIT:0] score_9_x26;
wire signed [DEBIT:0] score_9_x27;
wire signed [DEBIT:0] score_9_x28;
wire signed [DEBIT:0] score_9_x29;
wire signed [DEBIT:0] score_9_x30;
wire signed [DEBIT:0] score_9_x31;
wire signed [DEBIT:0] score_9_x32;
wire signed [DEBIT:0] score_9_x33;
wire signed [DEBIT:0] score_9_x34;
wire signed [DEBIT:0] score_9_x35;
wire signed [DEBIT:0] score_9_x36;
wire signed [DEBIT:0] score_9_x37;
wire signed [DEBIT:0] score_9_x38;
wire signed [DEBIT:0] score_9_x39;
wire signed [DEBIT:0] score_9_x40;
wire signed [DEBIT:0] score_9_x41;
wire signed [DEBIT:0] score_9_x42;
wire signed [DEBIT:0] score_9_x43;
wire signed [DEBIT:0] score_9_x44;
wire signed [DEBIT:0] score_9_x45;
wire signed [DEBIT:0] score_9_x46;
wire signed [DEBIT:0] score_9_x47;
wire signed [DEBIT:0] score_9_x48;
wire signed [DEBIT:0] score_9_x49;
wire signed [DEBIT:0] score_9_x50;
wire signed [DEBIT:0] score_9_x51;
wire signed [DEBIT:0] score_9_x52;
wire signed [DEBIT:0] score_9_x53;
wire signed [DEBIT:0] score_9_x54;
wire signed [DEBIT:0] score_9_x55;
wire signed [DEBIT:0] score_9_x56;
wire signed [DEBIT:0] score_9_x57;
wire signed [DEBIT:0] score_9_x58;
wire signed [DEBIT:0] score_9_x59;
wire signed [DEBIT:0] score_9_x60;
wire signed [DEBIT:0] score_9_x61;
wire signed [DEBIT:0] score_9_x62;
wire signed [DEBIT:0] score_9_x63;
wire signed [DEBIT:0] score_9_x64;
wire signed [DEBIT:0] score_9_x65;
wire signed [DEBIT:0] score_9_x66;
wire signed [DEBIT:0] score_9_x67;
wire signed [DEBIT:0] score_9_x68;
wire signed [DEBIT:0] score_9_x69;
wire signed [DEBIT:0] score_9_x70;
wire signed [DEBIT:0] score_9_x71;
wire signed [DEBIT:0] score_9_x72;
wire signed [DEBIT:0] score_9_x73;
wire signed [DEBIT:0] score_9_x74;
wire signed [DEBIT:0] score_9_x75;
wire signed [DEBIT:0] score_9_x76;
wire signed [DEBIT:0] score_9_x77;
wire signed [DEBIT:0] score_9_x78;
wire signed [DEBIT:0] score_9_x79;
wire signed [DEBIT:0] score_9_x80;
wire signed [DEBIT:0] score_9_x81;
wire signed [DEBIT:0] score_9_x82;
wire signed [DEBIT:0] score_9_x83;
wire signed [DEBIT:0] score_9_x84;
wire signed [DEBIT:0] score_9_x85;
wire signed [DEBIT:0] score_9_x86;
wire signed [DEBIT:0] score_9_x87;
wire signed [DEBIT:0] score_9_x88;
wire signed [DEBIT:0] score_9_x89;
wire signed [DEBIT:0] score_9_x90;
wire signed [DEBIT:0] score_9_x91;
wire signed [DEBIT:0] score_9_x92;
wire signed [DEBIT:0] score_9_x93;
wire signed [DEBIT:0] score_9_x94;
wire signed [DEBIT:0] score_9_x95;
wire signed [DEBIT:0] score_9_x96;
wire signed [DEBIT:0] score_9_x97;
wire signed [DEBIT:0] score_9_x98;
wire signed [DEBIT:0] score_9_x99;
wire signed [DEBIT:0] score_9_x100;
wire signed [DEBIT:0] score_9_x101;
wire signed [DEBIT:0] score_9_x102;
wire signed [DEBIT:0] score_9_x103;
wire signed [DEBIT:0] score_9_x104;
wire signed [DEBIT:0] score_9_x105;
wire signed [DEBIT:0] score_9_x106;
wire signed [DEBIT:0] score_9_x107;
wire signed [DEBIT:0] score_9_x108;
wire signed [DEBIT:0] score_9_x109;
wire signed [DEBIT:0] score_9_x110;
wire signed [DEBIT:0] score_9_x111;
wire signed [DEBIT:0] score_9_x112;
wire signed [DEBIT:0] score_9_x113;
wire signed [DEBIT:0] score_9_x114;
wire signed [DEBIT:0] score_9_x115;
wire signed [DEBIT:0] score_9_x116;
wire signed [DEBIT:0] score_9_x117;
wire signed [DEBIT:0] score_9_x118;
wire signed [DEBIT:0] score_9_x119;
wire signed [DEBIT:0] score_9_x120;
wire signed [DEBIT:0] score_9_x121;
wire signed [DEBIT:0] score_9_x122;
wire signed [DEBIT:0] score_9_x123;
wire signed [DEBIT:0] score_9_x124;
wire signed [DEBIT:0] score_9_x125;
wire signed [DEBIT:0] score_9_x126;
wire signed [DEBIT:0] score_9_x127;
wire signed [DEBIT:0] score_9_x128;
wire signed [DEBIT:0] score_9_x129;
wire signed [DEBIT:0] score_9_x130;
wire signed [DEBIT:0] score_9_x131;
wire signed [DEBIT:0] score_9_x132;
wire signed [DEBIT:0] score_9_x133;
wire signed [DEBIT:0] score_9_x134;
wire signed [DEBIT:0] score_9_x135;
wire signed [DEBIT:0] score_9_x136;
wire signed [DEBIT:0] score_9_x137;
wire signed [DEBIT:0] score_9_x138;
wire signed [DEBIT:0] score_9_x139;
wire signed [DEBIT:0] score_9_x140;
wire signed [DEBIT:0] score_9_x141;
wire signed [DEBIT:0] score_9_x142;
wire signed [DEBIT:0] score_9_x143;
wire signed [DEBIT:0] score_9_x144;
wire signed [DEBIT:0] score_9_x145;
wire signed [DEBIT:0] score_9_x146;
wire signed [DEBIT:0] score_9_x147;
wire signed [DEBIT:0] score_9_x148;
wire signed [DEBIT:0] score_9_x149;
wire signed [DEBIT:0] score_9_x150;
wire signed [DEBIT:0] score_9_x151;
wire signed [DEBIT:0] score_9_x152;
wire signed [DEBIT:0] score_9_x153;
wire signed [DEBIT:0] score_9_x154;
wire signed [DEBIT:0] score_9_x155;
wire signed [DEBIT:0] score_9_x156;
wire signed [DEBIT:0] score_9_x157;
wire signed [DEBIT:0] score_9_x158;
wire signed [DEBIT:0] score_9_x159;
wire signed [DEBIT:0] score_9_x160;
wire signed [DEBIT:0] score_9_x161;
wire signed [DEBIT:0] score_9_x162;
wire signed [DEBIT:0] score_9_x163;
wire signed [DEBIT:0] score_9_x164;
wire signed [DEBIT:0] score_9_x165;
wire signed [DEBIT:0] score_9_x166;
wire signed [DEBIT:0] score_9_x167;
wire signed [DEBIT:0] score_9_x168;
wire signed [DEBIT:0] score_9_x169;
wire signed [DEBIT:0] score_9_x170;
wire signed [DEBIT:0] score_9_x171;
wire signed [DEBIT:0] score_9_x172;
wire signed [DEBIT:0] score_9_x173;
wire signed [DEBIT:0] score_9_x174;
wire signed [DEBIT:0] score_9_x175;
wire signed [DEBIT:0] score_9_x176;
wire signed [DEBIT:0] score_9_x177;
wire signed [DEBIT:0] score_9_x178;
wire signed [DEBIT:0] score_9_x179;
wire signed [DEBIT:0] score_9_x180;
wire signed [DEBIT:0] score_9_x181;
wire signed [DEBIT:0] score_9_x182;
wire signed [DEBIT:0] score_9_x183;
wire signed [DEBIT:0] score_9_x184;
wire signed [DEBIT:0] score_9_x185;
wire signed [DEBIT:0] score_9_x186;
wire signed [DEBIT:0] score_9_x187;
wire signed [DEBIT:0] score_9_x188;
wire signed [DEBIT:0] score_9_x189;
wire signed [DEBIT:0] score_9_x190;
wire signed [DEBIT:0] score_9_x191;
wire signed [DEBIT:0] score_9_x192;
wire signed [DEBIT:0] score_9_x193;
wire signed [DEBIT:0] score_9_x194;
wire signed [DEBIT:0] score_9_x195;
wire signed [DEBIT:0] score_9_x196;
wire signed [DEBIT:0] score_9_x197;
wire signed [DEBIT:0] score_9_x198;
wire signed [DEBIT:0] score_9_x199;
wire signed [DEBIT:0] score_9_x200;
wire signed [DEBIT:0] score_9_x201;
wire signed [DEBIT:0] score_9_x202;
wire signed [DEBIT:0] score_9_x203;
wire signed [DEBIT:0] score_9_x204;
wire signed [DEBIT:0] score_9_x205;
wire signed [DEBIT:0] score_9_x206;
wire signed [DEBIT:0] score_9_x207;
wire signed [DEBIT:0] score_9_x208;
wire signed [DEBIT:0] score_9_x209;
wire signed [DEBIT:0] score_9_x210;
wire signed [DEBIT:0] score_9_x211;
wire signed [DEBIT:0] score_9_x212;
wire signed [DEBIT:0] score_9_x213;
wire signed [DEBIT:0] score_9_x214;
wire signed [DEBIT:0] score_9_x215;
wire signed [DEBIT:0] score_9_x216;
wire signed [DEBIT:0] score_9_x217;
wire signed [DEBIT:0] score_9_x218;
wire signed [DEBIT:0] score_9_x219;
wire signed [DEBIT:0] score_9_x220;
wire signed [DEBIT:0] score_9_x221;
wire signed [DEBIT:0] score_9_x222;
wire signed [DEBIT:0] score_9_x223;
wire signed [DEBIT:0] score_9_x224;
wire signed [DEBIT:0] score_9_x225;
wire signed [DEBIT:0] score_9_x226;
wire signed [DEBIT:0] score_9_x227;
wire signed [DEBIT:0] score_9_x228;
wire signed [DEBIT:0] score_9_x229;
wire signed [DEBIT:0] score_9_x230;
wire signed [DEBIT:0] score_9_x231;
wire signed [DEBIT:0] score_9_x232;
wire signed [DEBIT:0] score_9_x233;
wire signed [DEBIT:0] score_9_x234;
wire signed [DEBIT:0] score_9_x235;
wire signed [DEBIT:0] score_9_x236;
wire signed [DEBIT:0] score_9_x237;
wire signed [DEBIT:0] score_9_x238;
wire signed [DEBIT:0] score_9_x239;
wire signed [DEBIT:0] score_9_x240;
wire signed [DEBIT:0] score_9_x241;
wire signed [DEBIT:0] score_9_x242;
wire signed [DEBIT:0] score_9_x243;
wire signed [DEBIT:0] score_9_x244;
wire signed [DEBIT:0] score_9_x245;
wire signed [DEBIT:0] score_9_x246;
wire signed [DEBIT:0] score_9_x247;
wire signed [DEBIT:0] score_9_x248;
wire signed [DEBIT:0] score_9_x249;
wire signed [DEBIT:0] score_9_x250;
wire signed [DEBIT:0] score_9_x251;
wire signed [DEBIT:0] score_9_x252;
wire signed [DEBIT:0] score_9_x253;
wire signed [DEBIT:0] score_9_x254;
wire signed [DEBIT:0] score_9_x255;
wire signed [DEBIT:0] score_9_x256;
wire signed [DEBIT:0] score_9_x257;
wire signed [DEBIT:0] score_9_x258;
wire signed [DEBIT:0] score_9_x259;
wire signed [DEBIT:0] score_9_x260;
wire signed [DEBIT:0] score_9_x261;
wire signed [DEBIT:0] score_9_x262;
wire signed [DEBIT:0] score_9_x263;
wire signed [DEBIT:0] score_9_x264;
wire signed [DEBIT:0] score_9_x265;
wire signed [DEBIT:0] score_9_x266;
wire signed [DEBIT:0] score_9_x267;
wire signed [DEBIT:0] score_9_x268;
wire signed [DEBIT:0] score_9_x269;
wire signed [DEBIT:0] score_9_x270;
wire signed [DEBIT:0] score_9_x271;
wire signed [DEBIT:0] score_9_x272;
wire signed [DEBIT:0] score_9_x273;
wire signed [DEBIT:0] score_9_x274;
wire signed [DEBIT:0] score_9_x275;
wire signed [DEBIT:0] score_9_x276;
wire signed [DEBIT:0] score_9_x277;
wire signed [DEBIT:0] score_9_x278;
wire signed [DEBIT:0] score_9_x279;
wire signed [DEBIT:0] score_9_x280;
wire signed [DEBIT:0] score_9_x281;
wire signed [DEBIT:0] score_9_x282;
wire signed [DEBIT:0] score_9_x283;
wire signed [DEBIT:0] score_9_x284;
wire signed [DEBIT:0] score_9_x285;
wire signed [DEBIT:0] score_9_x286;
wire signed [DEBIT:0] score_9_x287;
wire signed [DEBIT:0] score_9_x288;
wire signed [DEBIT:0] score_9_x289;
wire signed [DEBIT:0] score_9_x290;
wire signed [DEBIT:0] score_9_x291;
wire signed [DEBIT:0] score_9_x292;
wire signed [DEBIT:0] score_9_x293;
wire signed [DEBIT:0] score_9_x294;
wire signed [DEBIT:0] score_9_x295;
wire signed [DEBIT:0] score_9_x296;
wire signed [DEBIT:0] score_9_x297;
wire signed [DEBIT:0] score_9_x298;
wire signed [DEBIT:0] score_9_x299;
wire signed [DEBIT:0] score_9_x300;
wire signed [DEBIT:0] score_9_x301;
wire signed [DEBIT:0] score_9_x302;
wire signed [DEBIT:0] score_9_x303;
wire signed [DEBIT:0] score_9_x304;
wire signed [DEBIT:0] score_9_x305;
wire signed [DEBIT:0] score_9_x306;
wire signed [DEBIT:0] score_9_x307;
wire signed [DEBIT:0] score_9_x308;
wire signed [DEBIT:0] score_9_x309;
wire signed [DEBIT:0] score_9_x310;
wire signed [DEBIT:0] score_9_x311;
wire signed [DEBIT:0] score_9_x312;
wire signed [DEBIT:0] score_9_x313;
wire signed [DEBIT:0] score_9_x314;
wire signed [DEBIT:0] score_9_x315;
wire signed [DEBIT:0] score_9_x316;
wire signed [DEBIT:0] score_9_x317;
wire signed [DEBIT:0] score_9_x318;
wire signed [DEBIT:0] score_9_x319;
wire signed [DEBIT:0] score_9_x320;
wire signed [DEBIT:0] score_9_x321;
wire signed [DEBIT:0] score_9_x322;
wire signed [DEBIT:0] score_9_x323;
wire signed [DEBIT:0] score_9_x324;
wire signed [DEBIT:0] score_9_x325;
wire signed [DEBIT:0] score_9_x326;
wire signed [DEBIT:0] score_9_x327;
wire signed [DEBIT:0] score_9_x328;
wire signed [DEBIT:0] score_9_x329;
wire signed [DEBIT:0] score_9_x330;
wire signed [DEBIT:0] score_9_x331;
wire signed [DEBIT:0] score_9_x332;
wire signed [DEBIT:0] score_9_x333;
wire signed [DEBIT:0] score_9_x334;
wire signed [DEBIT:0] score_9_x335;
wire signed [DEBIT:0] score_9_x336;
wire signed [DEBIT:0] score_9_x337;
wire signed [DEBIT:0] score_9_x338;
wire signed [DEBIT:0] score_9_x339;
wire signed [DEBIT:0] score_9_x340;
wire signed [DEBIT:0] score_9_x341;
wire signed [DEBIT:0] score_9_x342;
wire signed [DEBIT:0] score_9_x343;
wire signed [DEBIT:0] score_9_x344;
wire signed [DEBIT:0] score_9_x345;
wire signed [DEBIT:0] score_9_x346;
wire signed [DEBIT:0] score_9_x347;
wire signed [DEBIT:0] score_9_x348;
wire signed [DEBIT:0] score_9_x349;
wire signed [DEBIT:0] score_9_x350;
wire signed [DEBIT:0] score_9_x351;
wire signed [DEBIT:0] score_9_x352;
wire signed [DEBIT:0] score_9_x353;
wire signed [DEBIT:0] score_9_x354;
wire signed [DEBIT:0] score_9_x355;
wire signed [DEBIT:0] score_9_x356;
wire signed [DEBIT:0] score_9_x357;
wire signed [DEBIT:0] score_9_x358;
wire signed [DEBIT:0] score_9_x359;
wire signed [DEBIT:0] score_9_x360;
wire signed [DEBIT:0] score_9_x361;
wire signed [DEBIT:0] score_9_x362;
wire signed [DEBIT:0] score_9_x363;
wire signed [DEBIT:0] score_9_x364;
wire signed [DEBIT:0] score_9_x365;
wire signed [DEBIT:0] score_9_x366;
wire signed [DEBIT:0] score_9_x367;
wire signed [DEBIT:0] score_9_x368;
wire signed [DEBIT:0] score_9_x369;
wire signed [DEBIT:0] score_9_x370;
wire signed [DEBIT:0] score_9_x371;
wire signed [DEBIT:0] score_9_x372;
wire signed [DEBIT:0] score_9_x373;
wire signed [DEBIT:0] score_9_x374;
wire signed [DEBIT:0] score_9_x375;
wire signed [DEBIT:0] score_9_x376;
wire signed [DEBIT:0] score_9_x377;
wire signed [DEBIT:0] score_9_x378;
wire signed [DEBIT:0] score_9_x379;
wire signed [DEBIT:0] score_9_x380;
wire signed [DEBIT:0] score_9_x381;
wire signed [DEBIT:0] score_9_x382;
wire signed [DEBIT:0] score_9_x383;
wire signed [DEBIT:0] score_9_x384;
wire signed [DEBIT:0] score_9_x385;
wire signed [DEBIT:0] score_9_x386;
wire signed [DEBIT:0] score_9_x387;
wire signed [DEBIT:0] score_9_x388;
wire signed [DEBIT:0] score_9_x389;
wire signed [DEBIT:0] score_9_x390;
wire signed [DEBIT:0] score_9_x391;
wire signed [DEBIT:0] score_9_x392;
wire signed [DEBIT:0] score_9_x393;
wire signed [DEBIT:0] score_9_x394;
wire signed [DEBIT:0] score_9_x395;
wire signed [DEBIT:0] score_9_x396;
wire signed [DEBIT:0] score_9_x397;
wire signed [DEBIT:0] score_9_x398;
wire signed [DEBIT:0] score_9_x399;
wire signed [DEBIT:0] score_9_x400;
wire signed [DEBIT:0] score_9_x401;
wire signed [DEBIT:0] score_9_x402;
wire signed [DEBIT:0] score_9_x403;
wire signed [DEBIT:0] score_9_x404;
wire signed [DEBIT:0] score_9_x405;
wire signed [DEBIT:0] score_9_x406;
wire signed [DEBIT:0] score_9_x407;
wire signed [DEBIT:0] score_9_x408;
wire signed [DEBIT:0] score_9_x409;
wire signed [DEBIT:0] score_9_x410;
wire signed [DEBIT:0] score_9_x411;
wire signed [DEBIT:0] score_9_x412;
wire signed [DEBIT:0] score_9_x413;
wire signed [DEBIT:0] score_9_x414;
wire signed [DEBIT:0] score_9_x415;
wire signed [DEBIT:0] score_9_x416;
wire signed [DEBIT:0] score_9_x417;
wire signed [DEBIT:0] score_9_x418;
wire signed [DEBIT:0] score_9_x419;
wire signed [DEBIT:0] score_9_x420;
wire signed [DEBIT:0] score_9_x421;
wire signed [DEBIT:0] score_9_x422;
wire signed [DEBIT:0] score_9_x423;
wire signed [DEBIT:0] score_9_x424;
wire signed [DEBIT:0] score_9_x425;
wire signed [DEBIT:0] score_9_x426;
wire signed [DEBIT:0] score_9_x427;
wire signed [DEBIT:0] score_9_x428;
wire signed [DEBIT:0] score_9_x429;
wire signed [DEBIT:0] score_9_x430;
wire signed [DEBIT:0] score_9_x431;
wire signed [DEBIT:0] score_9_x432;
wire signed [DEBIT:0] score_9_x433;
wire signed [DEBIT:0] score_9_x434;
wire signed [DEBIT:0] score_9_x435;
wire signed [DEBIT:0] score_9_x436;
wire signed [DEBIT:0] score_9_x437;
wire signed [DEBIT:0] score_9_x438;
wire signed [DEBIT:0] score_9_x439;
wire signed [DEBIT:0] score_9_x440;
wire signed [DEBIT:0] score_9_x441;
wire signed [DEBIT:0] score_9_x442;
wire signed [DEBIT:0] score_9_x443;
wire signed [DEBIT:0] score_9_x444;
wire signed [DEBIT:0] score_9_x445;
wire signed [DEBIT:0] score_9_x446;
wire signed [DEBIT:0] score_9_x447;
wire signed [DEBIT:0] score_9_x448;
wire signed [DEBIT:0] score_9_x449;
wire signed [DEBIT:0] score_9_x450;
wire signed [DEBIT:0] score_9_x451;
wire signed [DEBIT:0] score_9_x452;
wire signed [DEBIT:0] score_9_x453;
wire signed [DEBIT:0] score_9_x454;
wire signed [DEBIT:0] score_9_x455;
wire signed [DEBIT:0] score_9_x456;
wire signed [DEBIT:0] score_9_x457;
wire signed [DEBIT:0] score_9_x458;
wire signed [DEBIT:0] score_9_x459;
wire signed [DEBIT:0] score_9_x460;
wire signed [DEBIT:0] score_9_x461;
wire signed [DEBIT:0] score_9_x462;
wire signed [DEBIT:0] score_9_x463;
wire signed [DEBIT:0] score_9_x464;
wire signed [DEBIT:0] score_9_x465;
wire signed [DEBIT:0] score_9_x466;
wire signed [DEBIT:0] score_9_x467;
wire signed [DEBIT:0] score_9_x468;
wire signed [DEBIT:0] score_9_x469;
wire signed [DEBIT:0] score_9_x470;
wire signed [DEBIT:0] score_9_x471;
wire signed [DEBIT:0] score_9_x472;
wire signed [DEBIT:0] score_9_x473;
wire signed [DEBIT:0] score_9_x474;
wire signed [DEBIT:0] score_9_x475;
wire signed [DEBIT:0] score_9_x476;
wire signed [DEBIT:0] score_9_x477;
wire signed [DEBIT:0] score_9_x478;
wire signed [DEBIT:0] score_9_x479;
wire signed [DEBIT:0] score_9_x480;
wire signed [DEBIT:0] score_9_x481;
wire signed [DEBIT:0] score_9_x482;
wire signed [DEBIT:0] score_9_x483;
wire signed [DEBIT:0] score_9_x484;
wire signed [DEBIT:0] score_9_x485;
wire signed [DEBIT:0] score_9_x486;
wire signed [DEBIT:0] score_9_x487;
wire signed [DEBIT:0] score_9_x488;
wire signed [DEBIT:0] score_9_x489;
wire signed [DEBIT:0] score_9_x490;
wire signed [DEBIT:0] score_9_x491;
wire signed [DEBIT:0] score_9_x492;
wire signed [DEBIT:0] score_9_x493;
wire signed [DEBIT:0] score_9_x494;
wire signed [DEBIT:0] score_9_x495;
wire signed [DEBIT:0] score_9_x496;
wire signed [DEBIT:0] score_9_x497;
wire signed [DEBIT:0] score_9_x498;
wire signed [DEBIT:0] score_9_x499;
wire signed [DEBIT:0] score_9_x500;
wire signed [DEBIT:0] score_9_x501;
wire signed [DEBIT:0] score_9_x502;
wire signed [DEBIT:0] score_9_x503;
wire signed [DEBIT:0] score_9_x504;
wire signed [DEBIT:0] score_9_x505;
wire signed [DEBIT:0] score_9_x506;
wire signed [DEBIT:0] score_9_x507;
wire signed [DEBIT:0] score_9_x508;
wire signed [DEBIT:0] score_9_x509;
wire signed [DEBIT:0] score_9_x510;
wire signed [DEBIT:0] score_9_x511;
wire signed [DEBIT:0] score_9_x512;
wire signed [DEBIT:0] score_9_x513;
wire signed [DEBIT:0] score_9_x514;
wire signed [DEBIT:0] score_9_x515;
wire signed [DEBIT:0] score_9_x516;
wire signed [DEBIT:0] score_9_x517;
wire signed [DEBIT:0] score_9_x518;
wire signed [DEBIT:0] score_9_x519;
wire signed [DEBIT:0] score_9_x520;
wire signed [DEBIT:0] score_9_x521;
wire signed [DEBIT:0] score_9_x522;
wire signed [DEBIT:0] score_9_x523;
wire signed [DEBIT:0] score_9_x524;
wire signed [DEBIT:0] score_9_x525;
wire signed [DEBIT:0] score_9_x526;
wire signed [DEBIT:0] score_9_x527;
wire signed [DEBIT:0] score_9_x528;
wire signed [DEBIT:0] score_9_x529;
wire signed [DEBIT:0] score_9_x530;
wire signed [DEBIT:0] score_9_x531;
wire signed [DEBIT:0] score_9_x532;
wire signed [DEBIT:0] score_9_x533;
wire signed [DEBIT:0] score_9_x534;
wire signed [DEBIT:0] score_9_x535;
wire signed [DEBIT:0] score_9_x536;
wire signed [DEBIT:0] score_9_x537;
wire signed [DEBIT:0] score_9_x538;
wire signed [DEBIT:0] score_9_x539;
wire signed [DEBIT:0] score_9_x540;
wire signed [DEBIT:0] score_9_x541;
wire signed [DEBIT:0] score_9_x542;
wire signed [DEBIT:0] score_9_x543;
wire signed [DEBIT:0] score_9_x544;
wire signed [DEBIT:0] score_9_x545;
wire signed [DEBIT:0] score_9_x546;
wire signed [DEBIT:0] score_9_x547;
wire signed [DEBIT:0] score_9_x548;
wire signed [DEBIT:0] score_9_x549;
wire signed [DEBIT:0] score_9_x550;
wire signed [DEBIT:0] score_9_x551;
wire signed [DEBIT:0] score_9_x552;
wire signed [DEBIT:0] score_9_x553;
wire signed [DEBIT:0] score_9_x554;
wire signed [DEBIT:0] score_9_x555;
wire signed [DEBIT:0] score_9_x556;
wire signed [DEBIT:0] score_9_x557;
wire signed [DEBIT:0] score_9_x558;
wire signed [DEBIT:0] score_9_x559;
wire signed [DEBIT:0] score_9_x560;
wire signed [DEBIT:0] score_9_x561;
wire signed [DEBIT:0] score_9_x562;
wire signed [DEBIT:0] score_9_x563;
wire signed [DEBIT:0] score_9_x564;
wire signed [DEBIT:0] score_9_x565;
wire signed [DEBIT:0] score_9_x566;
wire signed [DEBIT:0] score_9_x567;
wire signed [DEBIT:0] score_9_x568;
wire signed [DEBIT:0] score_9_x569;
wire signed [DEBIT:0] score_9_x570;
wire signed [DEBIT:0] score_9_x571;
wire signed [DEBIT:0] score_9_x572;
wire signed [DEBIT:0] score_9_x573;
wire signed [DEBIT:0] score_9_x574;
wire signed [DEBIT:0] score_9_x575;
wire signed [DEBIT:0] score_9_x576;
wire signed [DEBIT:0] score_9_x577;
wire signed [DEBIT:0] score_9_x578;
wire signed [DEBIT:0] score_9_x579;
wire signed [DEBIT:0] score_9_x580;
wire signed [DEBIT:0] score_9_x581;
wire signed [DEBIT:0] score_9_x582;
wire signed [DEBIT:0] score_9_x583;
wire signed [DEBIT:0] score_9_x584;
wire signed [DEBIT:0] score_9_x585;
wire signed [DEBIT:0] score_9_x586;
wire signed [DEBIT:0] score_9_x587;
wire signed [DEBIT:0] score_9_x588;
wire signed [DEBIT:0] score_9_x589;
wire signed [DEBIT:0] score_9_x590;
wire signed [DEBIT:0] score_9_x591;
wire signed [DEBIT:0] score_9_x592;
wire signed [DEBIT:0] score_9_x593;
wire signed [DEBIT:0] score_9_x594;
wire signed [DEBIT:0] score_9_x595;
wire signed [DEBIT:0] score_9_x596;
wire signed [DEBIT:0] score_9_x597;
wire signed [DEBIT:0] score_9_x598;
wire signed [DEBIT:0] score_9_x599;
wire signed [DEBIT:0] score_9_x600;
wire signed [DEBIT:0] score_9_x601;
wire signed [DEBIT:0] score_9_x602;
wire signed [DEBIT:0] score_9_x603;
wire signed [DEBIT:0] score_9_x604;
wire signed [DEBIT:0] score_9_x605;
wire signed [DEBIT:0] score_9_x606;
wire signed [DEBIT:0] score_9_x607;
wire signed [DEBIT:0] score_9_x608;
wire signed [DEBIT:0] score_9_x609;
wire signed [DEBIT:0] score_9_x610;
wire signed [DEBIT:0] score_9_x611;
wire signed [DEBIT:0] score_9_x612;
wire signed [DEBIT:0] score_9_x613;
wire signed [DEBIT:0] score_9_x614;
wire signed [DEBIT:0] score_9_x615;
wire signed [DEBIT:0] score_9_x616;
wire signed [DEBIT:0] score_9_x617;
wire signed [DEBIT:0] score_9_x618;
wire signed [DEBIT:0] score_9_x619;
wire signed [DEBIT:0] score_9_x620;
wire signed [DEBIT:0] score_9_x621;
wire signed [DEBIT:0] score_9_x622;
wire signed [DEBIT:0] score_9_x623;
wire signed [DEBIT:0] score_9_x624;
wire signed [DEBIT:0] score_9_x625;
wire signed [DEBIT:0] score_9_x626;
wire signed [DEBIT:0] score_9_x627;
wire signed [DEBIT:0] score_9_x628;
wire signed [DEBIT:0] score_9_x629;
wire signed [DEBIT:0] score_9_x630;
wire signed [DEBIT:0] score_9_x631;
wire signed [DEBIT:0] score_9_x632;
wire signed [DEBIT:0] score_9_x633;
wire signed [DEBIT:0] score_9_x634;
wire signed [DEBIT:0] score_9_x635;
wire signed [DEBIT:0] score_9_x636;
wire signed [DEBIT:0] score_9_x637;
wire signed [DEBIT:0] score_9_x638;
wire signed [DEBIT:0] score_9_x639;
wire signed [DEBIT:0] score_9_x640;
wire signed [DEBIT:0] score_9_x641;
wire signed [DEBIT:0] score_9_x642;
wire signed [DEBIT:0] score_9_x643;
wire signed [DEBIT:0] score_9_x644;
wire signed [DEBIT:0] score_9_x645;
wire signed [DEBIT:0] score_9_x646;
wire signed [DEBIT:0] score_9_x647;
wire signed [DEBIT:0] score_9_x648;
wire signed [DEBIT:0] score_9_x649;
wire signed [DEBIT:0] score_9_x650;
wire signed [DEBIT:0] score_9_x651;
wire signed [DEBIT:0] score_9_x652;
wire signed [DEBIT:0] score_9_x653;
wire signed [DEBIT:0] score_9_x654;
wire signed [DEBIT:0] score_9_x655;
wire signed [DEBIT:0] score_9_x656;
wire signed [DEBIT:0] score_9_x657;
wire signed [DEBIT:0] score_9_x658;
wire signed [DEBIT:0] score_9_x659;
wire signed [DEBIT:0] score_9_x660;
wire signed [DEBIT:0] score_9_x661;
wire signed [DEBIT:0] score_9_x662;
wire signed [DEBIT:0] score_9_x663;
wire signed [DEBIT:0] score_9_x664;
wire signed [DEBIT:0] score_9_x665;
wire signed [DEBIT:0] score_9_x666;
wire signed [DEBIT:0] score_9_x667;
wire signed [DEBIT:0] score_9_x668;
wire signed [DEBIT:0] score_9_x669;
wire signed [DEBIT:0] score_9_x670;
wire signed [DEBIT:0] score_9_x671;
wire signed [DEBIT:0] score_9_x672;
wire signed [DEBIT:0] score_9_x673;
wire signed [DEBIT:0] score_9_x674;
wire signed [DEBIT:0] score_9_x675;
wire signed [DEBIT:0] score_9_x676;
wire signed [DEBIT:0] score_9_x677;
wire signed [DEBIT:0] score_9_x678;
wire signed [DEBIT:0] score_9_x679;
wire signed [DEBIT:0] score_9_x680;
wire signed [DEBIT:0] score_9_x681;
wire signed [DEBIT:0] score_9_x682;
wire signed [DEBIT:0] score_9_x683;
wire signed [DEBIT:0] score_9_x684;
wire signed [DEBIT:0] score_9_x685;
wire signed [DEBIT:0] score_9_x686;
wire signed [DEBIT:0] score_9_x687;
wire signed [DEBIT:0] score_9_x688;
wire signed [DEBIT:0] score_9_x689;
wire signed [DEBIT:0] score_9_x690;
wire signed [DEBIT:0] score_9_x691;
wire signed [DEBIT:0] score_9_x692;
wire signed [DEBIT:0] score_9_x693;
wire signed [DEBIT:0] score_9_x694;
wire signed [DEBIT:0] score_9_x695;
wire signed [DEBIT:0] score_9_x696;
wire signed [DEBIT:0] score_9_x697;
wire signed [DEBIT:0] score_9_x698;
wire signed [DEBIT:0] score_9_x699;
wire signed [DEBIT:0] score_9_x700;
wire signed [DEBIT:0] score_9_x701;
wire signed [DEBIT:0] score_9_x702;
wire signed [DEBIT:0] score_9_x703;
wire signed [DEBIT:0] score_9_x704;
wire signed [DEBIT:0] score_9_x705;
wire signed [DEBIT:0] score_9_x706;
wire signed [DEBIT:0] score_9_x707;
wire signed [DEBIT:0] score_9_x708;
wire signed [DEBIT:0] score_9_x709;
wire signed [DEBIT:0] score_9_x710;
wire signed [DEBIT:0] score_9_x711;
wire signed [DEBIT:0] score_9_x712;
wire signed [DEBIT:0] score_9_x713;
wire signed [DEBIT:0] score_9_x714;
wire signed [DEBIT:0] score_9_x715;
wire signed [DEBIT:0] score_9_x716;
wire signed [DEBIT:0] score_9_x717;
wire signed [DEBIT:0] score_9_x718;
wire signed [DEBIT:0] score_9_x719;
wire signed [DEBIT:0] score_9_x720;
wire signed [DEBIT:0] score_9_x721;
wire signed [DEBIT:0] score_9_x722;
wire signed [DEBIT:0] score_9_x723;
wire signed [DEBIT:0] score_9_x724;
wire signed [DEBIT:0] score_9_x725;
wire signed [DEBIT:0] score_9_x726;
wire signed [DEBIT:0] score_9_x727;
wire signed [DEBIT:0] score_9_x728;
wire signed [DEBIT:0] score_9_x729;
wire signed [DEBIT:0] score_9_x730;
wire signed [DEBIT:0] score_9_x731;
wire signed [DEBIT:0] score_9_x732;
wire signed [DEBIT:0] score_9_x733;
wire signed [DEBIT:0] score_9_x734;
wire signed [DEBIT:0] score_9_x735;
wire signed [DEBIT:0] score_9_x736;
wire signed [DEBIT:0] score_9_x737;
wire signed [DEBIT:0] score_9_x738;
wire signed [DEBIT:0] score_9_x739;
wire signed [DEBIT:0] score_9_x740;
wire signed [DEBIT:0] score_9_x741;
wire signed [DEBIT:0] score_9_x742;
wire signed [DEBIT:0] score_9_x743;
wire signed [DEBIT:0] score_9_x744;
wire signed [DEBIT:0] score_9_x745;
wire signed [DEBIT:0] score_9_x746;
wire signed [DEBIT:0] score_9_x747;
wire signed [DEBIT:0] score_9_x748;
wire signed [DEBIT:0] score_9_x749;
wire signed [DEBIT:0] score_9_x750;
wire signed [DEBIT:0] score_9_x751;
wire signed [DEBIT:0] score_9_x752;
wire signed [DEBIT:0] score_9_x753;
wire signed [DEBIT:0] score_9_x754;
wire signed [DEBIT:0] score_9_x755;
wire signed [DEBIT:0] score_9_x756;
wire signed [DEBIT:0] score_9_x757;
wire signed [DEBIT:0] score_9_x758;
wire signed [DEBIT:0] score_9_x759;
wire signed [DEBIT:0] score_9_x760;
wire signed [DEBIT:0] score_9_x761;
wire signed [DEBIT:0] score_9_x762;
wire signed [DEBIT:0] score_9_x763;
wire signed [DEBIT:0] score_9_x764;
wire signed [DEBIT:0] score_9_x765;
wire signed [DEBIT:0] score_9_x766;
wire signed [DEBIT:0] score_9_x767;
wire signed [DEBIT:0] score_9_x768;
wire signed [DEBIT:0] score_9_x769;
wire signed [DEBIT:0] score_9_x770;
wire signed [DEBIT:0] score_9_x771;
wire signed [DEBIT:0] score_9_x772;
wire signed [DEBIT:0] score_9_x773;
wire signed [DEBIT:0] score_9_x774;
wire signed [DEBIT:0] score_9_x775;
wire signed [DEBIT:0] score_9_x776;
wire signed [DEBIT:0] score_9_x777;
wire signed [DEBIT:0] score_9_x778;
wire signed [DEBIT:0] score_9_x779;
wire signed [DEBIT:0] score_9_x780;
wire signed [DEBIT:0] score_9_x781;
wire signed [DEBIT:0] score_9_x782;
wire signed [DEBIT:0] score_9_x783;
wire signed [DEBIT:0] score_9_x784;

//=============================================================================
//****************************     Main Code    *******************************
//=============================================================================



//****************************    存入判断值    *******************************








always @ (posedge clk) begin
	if(rst_valid) begin
      res_0_sum <= 1'b0;
      res_1_sum <= 1'b0;
      res_2_sum <= 1'b0;
      res_3_sum <= 1'b0;
      res_4_sum <= 1'b0;
      res_5_sum <= 1'b0;
      res_6_sum <= 1'b0;
      res_7_sum <= 1'b0;
      res_8_sum <= 1'b0;
      res_9_sum <= 1'b0;
	end	
	else if(res_done_x1) begin
      res_0_sum <= res_0_sum + score_0_x1;
      res_1_sum <= res_1_sum + score_1_x1;
      res_2_sum <= res_2_sum + score_2_x1;
      res_3_sum <= res_3_sum + score_3_x1;
      res_4_sum <= res_4_sum + score_4_x1;
      res_5_sum <= res_5_sum + score_5_x1;
      res_6_sum <= res_6_sum + score_6_x1;
      res_7_sum <= res_7_sum + score_7_x1;
      res_8_sum <= res_8_sum + score_8_x1;
      res_9_sum <= res_9_sum + score_9_x1;
   end
   else if(res_done_x2) begin
      res_0_sum <= res_0_sum + score_0_x2;
      res_1_sum <= res_1_sum + score_1_x2;
      res_2_sum <= res_2_sum + score_2_x2;
      res_3_sum <= res_3_sum + score_3_x2;
      res_4_sum <= res_4_sum + score_4_x2;
      res_5_sum <= res_5_sum + score_5_x2;
      res_6_sum <= res_6_sum + score_6_x2;
      res_7_sum <= res_7_sum + score_7_x2;
      res_8_sum <= res_8_sum + score_8_x2;
      res_9_sum <= res_9_sum + score_9_x2;
   end
   else if(res_done_x3) begin
      res_0_sum <= res_0_sum + score_0_x3;
      res_1_sum <= res_1_sum + score_1_x3;
      res_2_sum <= res_2_sum + score_2_x3;
      res_3_sum <= res_3_sum + score_3_x3;
      res_4_sum <= res_4_sum + score_4_x3;
      res_5_sum <= res_5_sum + score_5_x3;
      res_6_sum <= res_6_sum + score_6_x3;
      res_7_sum <= res_7_sum + score_7_x3;
      res_8_sum <= res_8_sum + score_8_x3;
      res_9_sum <= res_9_sum + score_9_x3;
   end
   else if(res_done_x4) begin
      res_0_sum <= res_0_sum + score_0_x4;
      res_1_sum <= res_1_sum + score_1_x4;
      res_2_sum <= res_2_sum + score_2_x4;
      res_3_sum <= res_3_sum + score_3_x4;
      res_4_sum <= res_4_sum + score_4_x4;
      res_5_sum <= res_5_sum + score_5_x4;
      res_6_sum <= res_6_sum + score_6_x4;
      res_7_sum <= res_7_sum + score_7_x4;
      res_8_sum <= res_8_sum + score_8_x4;
      res_9_sum <= res_9_sum + score_9_x4;
   end
   else if(res_done_x5) begin
      res_0_sum <= res_0_sum + score_0_x5;
      res_1_sum <= res_1_sum + score_1_x5;
      res_2_sum <= res_2_sum + score_2_x5;
      res_3_sum <= res_3_sum + score_3_x5;
      res_4_sum <= res_4_sum + score_4_x5;
      res_5_sum <= res_5_sum + score_5_x5;
      res_6_sum <= res_6_sum + score_6_x5;
      res_7_sum <= res_7_sum + score_7_x5;
      res_8_sum <= res_8_sum + score_8_x5;
      res_9_sum <= res_9_sum + score_9_x5;
   end
   else if(res_done_x6) begin
      res_0_sum <= res_0_sum + score_0_x6;
      res_1_sum <= res_1_sum + score_1_x6;
      res_2_sum <= res_2_sum + score_2_x6;
      res_3_sum <= res_3_sum + score_3_x6;
      res_4_sum <= res_4_sum + score_4_x6;
      res_5_sum <= res_5_sum + score_5_x6;
      res_6_sum <= res_6_sum + score_6_x6;
      res_7_sum <= res_7_sum + score_7_x6;
      res_8_sum <= res_8_sum + score_8_x6;
      res_9_sum <= res_9_sum + score_9_x6;
   end
   else if(res_done_x7) begin
      res_0_sum <= res_0_sum + score_0_x7;
      res_1_sum <= res_1_sum + score_1_x7;
      res_2_sum <= res_2_sum + score_2_x7;
      res_3_sum <= res_3_sum + score_3_x7;
      res_4_sum <= res_4_sum + score_4_x7;
      res_5_sum <= res_5_sum + score_5_x7;
      res_6_sum <= res_6_sum + score_6_x7;
      res_7_sum <= res_7_sum + score_7_x7;
      res_8_sum <= res_8_sum + score_8_x7;
      res_9_sum <= res_9_sum + score_9_x7;
   end
   else if(res_done_x8) begin
      res_0_sum <= res_0_sum + score_0_x8;
      res_1_sum <= res_1_sum + score_1_x8;
      res_2_sum <= res_2_sum + score_2_x8;
      res_3_sum <= res_3_sum + score_3_x8;
      res_4_sum <= res_4_sum + score_4_x8;
      res_5_sum <= res_5_sum + score_5_x8;
      res_6_sum <= res_6_sum + score_6_x8;
      res_7_sum <= res_7_sum + score_7_x8;
      res_8_sum <= res_8_sum + score_8_x8;
      res_9_sum <= res_9_sum + score_9_x8;
   end
   else if(res_done_x9) begin
      res_0_sum <= res_0_sum + score_0_x9;
      res_1_sum <= res_1_sum + score_1_x9;
      res_2_sum <= res_2_sum + score_2_x9;
      res_3_sum <= res_3_sum + score_3_x9;
      res_4_sum <= res_4_sum + score_4_x9;
      res_5_sum <= res_5_sum + score_5_x9;
      res_6_sum <= res_6_sum + score_6_x9;
      res_7_sum <= res_7_sum + score_7_x9;
      res_8_sum <= res_8_sum + score_8_x9;
      res_9_sum <= res_9_sum + score_9_x9;
   end
   else if(res_done_x10) begin
      res_0_sum <= res_0_sum + score_0_x10;
      res_1_sum <= res_1_sum + score_1_x10;
      res_2_sum <= res_2_sum + score_2_x10;
      res_3_sum <= res_3_sum + score_3_x10;
      res_4_sum <= res_4_sum + score_4_x10;
      res_5_sum <= res_5_sum + score_5_x10;
      res_6_sum <= res_6_sum + score_6_x10;
      res_7_sum <= res_7_sum + score_7_x10;
      res_8_sum <= res_8_sum + score_8_x10;
      res_9_sum <= res_9_sum + score_9_x10;
   end
   else if(res_done_x11) begin
      res_0_sum <= res_0_sum + score_0_x11;
      res_1_sum <= res_1_sum + score_1_x11;
      res_2_sum <= res_2_sum + score_2_x11;
      res_3_sum <= res_3_sum + score_3_x11;
      res_4_sum <= res_4_sum + score_4_x11;
      res_5_sum <= res_5_sum + score_5_x11;
      res_6_sum <= res_6_sum + score_6_x11;
      res_7_sum <= res_7_sum + score_7_x11;
      res_8_sum <= res_8_sum + score_8_x11;
      res_9_sum <= res_9_sum + score_9_x11;
   end
   else if(res_done_x12) begin
      res_0_sum <= res_0_sum + score_0_x12;
      res_1_sum <= res_1_sum + score_1_x12;
      res_2_sum <= res_2_sum + score_2_x12;
      res_3_sum <= res_3_sum + score_3_x12;
      res_4_sum <= res_4_sum + score_4_x12;
      res_5_sum <= res_5_sum + score_5_x12;
      res_6_sum <= res_6_sum + score_6_x12;
      res_7_sum <= res_7_sum + score_7_x12;
      res_8_sum <= res_8_sum + score_8_x12;
      res_9_sum <= res_9_sum + score_9_x12;
   end
   else if(res_done_x13) begin
      res_0_sum <= res_0_sum + score_0_x13;
      res_1_sum <= res_1_sum + score_1_x13;
      res_2_sum <= res_2_sum + score_2_x13;
      res_3_sum <= res_3_sum + score_3_x13;
      res_4_sum <= res_4_sum + score_4_x13;
      res_5_sum <= res_5_sum + score_5_x13;
      res_6_sum <= res_6_sum + score_6_x13;
      res_7_sum <= res_7_sum + score_7_x13;
      res_8_sum <= res_8_sum + score_8_x13;
      res_9_sum <= res_9_sum + score_9_x13;
   end
   else if(res_done_x14) begin
      res_0_sum <= res_0_sum + score_0_x14;
      res_1_sum <= res_1_sum + score_1_x14;
      res_2_sum <= res_2_sum + score_2_x14;
      res_3_sum <= res_3_sum + score_3_x14;
      res_4_sum <= res_4_sum + score_4_x14;
      res_5_sum <= res_5_sum + score_5_x14;
      res_6_sum <= res_6_sum + score_6_x14;
      res_7_sum <= res_7_sum + score_7_x14;
      res_8_sum <= res_8_sum + score_8_x14;
      res_9_sum <= res_9_sum + score_9_x14;
   end
   else if(res_done_x15) begin
      res_0_sum <= res_0_sum + score_0_x15;
      res_1_sum <= res_1_sum + score_1_x15;
      res_2_sum <= res_2_sum + score_2_x15;
      res_3_sum <= res_3_sum + score_3_x15;
      res_4_sum <= res_4_sum + score_4_x15;
      res_5_sum <= res_5_sum + score_5_x15;
      res_6_sum <= res_6_sum + score_6_x15;
      res_7_sum <= res_7_sum + score_7_x15;
      res_8_sum <= res_8_sum + score_8_x15;
      res_9_sum <= res_9_sum + score_9_x15;
   end
   else if(res_done_x16) begin
      res_0_sum <= res_0_sum + score_0_x16;
      res_1_sum <= res_1_sum + score_1_x16;
      res_2_sum <= res_2_sum + score_2_x16;
      res_3_sum <= res_3_sum + score_3_x16;
      res_4_sum <= res_4_sum + score_4_x16;
      res_5_sum <= res_5_sum + score_5_x16;
      res_6_sum <= res_6_sum + score_6_x16;
      res_7_sum <= res_7_sum + score_7_x16;
      res_8_sum <= res_8_sum + score_8_x16;
      res_9_sum <= res_9_sum + score_9_x16;
   end
   else if(res_done_x17) begin
      res_0_sum <= res_0_sum + score_0_x17;
      res_1_sum <= res_1_sum + score_1_x17;
      res_2_sum <= res_2_sum + score_2_x17;
      res_3_sum <= res_3_sum + score_3_x17;
      res_4_sum <= res_4_sum + score_4_x17;
      res_5_sum <= res_5_sum + score_5_x17;
      res_6_sum <= res_6_sum + score_6_x17;
      res_7_sum <= res_7_sum + score_7_x17;
      res_8_sum <= res_8_sum + score_8_x17;
      res_9_sum <= res_9_sum + score_9_x17;
   end
   else if(res_done_x18) begin
      res_0_sum <= res_0_sum + score_0_x18;
      res_1_sum <= res_1_sum + score_1_x18;
      res_2_sum <= res_2_sum + score_2_x18;
      res_3_sum <= res_3_sum + score_3_x18;
      res_4_sum <= res_4_sum + score_4_x18;
      res_5_sum <= res_5_sum + score_5_x18;
      res_6_sum <= res_6_sum + score_6_x18;
      res_7_sum <= res_7_sum + score_7_x18;
      res_8_sum <= res_8_sum + score_8_x18;
      res_9_sum <= res_9_sum + score_9_x18;
   end
   else if(res_done_x19) begin
      res_0_sum <= res_0_sum + score_0_x19;
      res_1_sum <= res_1_sum + score_1_x19;
      res_2_sum <= res_2_sum + score_2_x19;
      res_3_sum <= res_3_sum + score_3_x19;
      res_4_sum <= res_4_sum + score_4_x19;
      res_5_sum <= res_5_sum + score_5_x19;
      res_6_sum <= res_6_sum + score_6_x19;
      res_7_sum <= res_7_sum + score_7_x19;
      res_8_sum <= res_8_sum + score_8_x19;
      res_9_sum <= res_9_sum + score_9_x19;
   end
   else if(res_done_x20) begin
      res_0_sum <= res_0_sum + score_0_x20;
      res_1_sum <= res_1_sum + score_1_x20;
      res_2_sum <= res_2_sum + score_2_x20;
      res_3_sum <= res_3_sum + score_3_x20;
      res_4_sum <= res_4_sum + score_4_x20;
      res_5_sum <= res_5_sum + score_5_x20;
      res_6_sum <= res_6_sum + score_6_x20;
      res_7_sum <= res_7_sum + score_7_x20;
      res_8_sum <= res_8_sum + score_8_x20;
      res_9_sum <= res_9_sum + score_9_x20;
   end
   else if(res_done_x21) begin
      res_0_sum <= res_0_sum + score_0_x21;
      res_1_sum <= res_1_sum + score_1_x21;
      res_2_sum <= res_2_sum + score_2_x21;
      res_3_sum <= res_3_sum + score_3_x21;
      res_4_sum <= res_4_sum + score_4_x21;
      res_5_sum <= res_5_sum + score_5_x21;
      res_6_sum <= res_6_sum + score_6_x21;
      res_7_sum <= res_7_sum + score_7_x21;
      res_8_sum <= res_8_sum + score_8_x21;
      res_9_sum <= res_9_sum + score_9_x21;
   end
   else if(res_done_x22) begin
      res_0_sum <= res_0_sum + score_0_x22;
      res_1_sum <= res_1_sum + score_1_x22;
      res_2_sum <= res_2_sum + score_2_x22;
      res_3_sum <= res_3_sum + score_3_x22;
      res_4_sum <= res_4_sum + score_4_x22;
      res_5_sum <= res_5_sum + score_5_x22;
      res_6_sum <= res_6_sum + score_6_x22;
      res_7_sum <= res_7_sum + score_7_x22;
      res_8_sum <= res_8_sum + score_8_x22;
      res_9_sum <= res_9_sum + score_9_x22;
   end
   else if(res_done_x23) begin
      res_0_sum <= res_0_sum + score_0_x23;
      res_1_sum <= res_1_sum + score_1_x23;
      res_2_sum <= res_2_sum + score_2_x23;
      res_3_sum <= res_3_sum + score_3_x23;
      res_4_sum <= res_4_sum + score_4_x23;
      res_5_sum <= res_5_sum + score_5_x23;
      res_6_sum <= res_6_sum + score_6_x23;
      res_7_sum <= res_7_sum + score_7_x23;
      res_8_sum <= res_8_sum + score_8_x23;
      res_9_sum <= res_9_sum + score_9_x23;
   end
   else if(res_done_x24) begin
      res_0_sum <= res_0_sum + score_0_x24;
      res_1_sum <= res_1_sum + score_1_x24;
      res_2_sum <= res_2_sum + score_2_x24;
      res_3_sum <= res_3_sum + score_3_x24;
      res_4_sum <= res_4_sum + score_4_x24;
      res_5_sum <= res_5_sum + score_5_x24;
      res_6_sum <= res_6_sum + score_6_x24;
      res_7_sum <= res_7_sum + score_7_x24;
      res_8_sum <= res_8_sum + score_8_x24;
      res_9_sum <= res_9_sum + score_9_x24;
   end
   else if(res_done_x25) begin
      res_0_sum <= res_0_sum + score_0_x25;
      res_1_sum <= res_1_sum + score_1_x25;
      res_2_sum <= res_2_sum + score_2_x25;
      res_3_sum <= res_3_sum + score_3_x25;
      res_4_sum <= res_4_sum + score_4_x25;
      res_5_sum <= res_5_sum + score_5_x25;
      res_6_sum <= res_6_sum + score_6_x25;
      res_7_sum <= res_7_sum + score_7_x25;
      res_8_sum <= res_8_sum + score_8_x25;
      res_9_sum <= res_9_sum + score_9_x25;
   end
   else if(res_done_x26) begin
      res_0_sum <= res_0_sum + score_0_x26;
      res_1_sum <= res_1_sum + score_1_x26;
      res_2_sum <= res_2_sum + score_2_x26;
      res_3_sum <= res_3_sum + score_3_x26;
      res_4_sum <= res_4_sum + score_4_x26;
      res_5_sum <= res_5_sum + score_5_x26;
      res_6_sum <= res_6_sum + score_6_x26;
      res_7_sum <= res_7_sum + score_7_x26;
      res_8_sum <= res_8_sum + score_8_x26;
      res_9_sum <= res_9_sum + score_9_x26;
   end
   else if(res_done_x27) begin
      res_0_sum <= res_0_sum + score_0_x27;
      res_1_sum <= res_1_sum + score_1_x27;
      res_2_sum <= res_2_sum + score_2_x27;
      res_3_sum <= res_3_sum + score_3_x27;
      res_4_sum <= res_4_sum + score_4_x27;
      res_5_sum <= res_5_sum + score_5_x27;
      res_6_sum <= res_6_sum + score_6_x27;
      res_7_sum <= res_7_sum + score_7_x27;
      res_8_sum <= res_8_sum + score_8_x27;
      res_9_sum <= res_9_sum + score_9_x27;
   end
   else if(res_done_x28) begin
      res_0_sum <= res_0_sum + score_0_x28;
      res_1_sum <= res_1_sum + score_1_x28;
      res_2_sum <= res_2_sum + score_2_x28;
      res_3_sum <= res_3_sum + score_3_x28;
      res_4_sum <= res_4_sum + score_4_x28;
      res_5_sum <= res_5_sum + score_5_x28;
      res_6_sum <= res_6_sum + score_6_x28;
      res_7_sum <= res_7_sum + score_7_x28;
      res_8_sum <= res_8_sum + score_8_x28;
      res_9_sum <= res_9_sum + score_9_x28;
   end
   else if(res_done_x29) begin
      res_0_sum <= res_0_sum + score_0_x29;
      res_1_sum <= res_1_sum + score_1_x29;
      res_2_sum <= res_2_sum + score_2_x29;
      res_3_sum <= res_3_sum + score_3_x29;
      res_4_sum <= res_4_sum + score_4_x29;
      res_5_sum <= res_5_sum + score_5_x29;
      res_6_sum <= res_6_sum + score_6_x29;
      res_7_sum <= res_7_sum + score_7_x29;
      res_8_sum <= res_8_sum + score_8_x29;
      res_9_sum <= res_9_sum + score_9_x29;
   end
   else if(res_done_x30) begin
      res_0_sum <= res_0_sum + score_0_x30;
      res_1_sum <= res_1_sum + score_1_x30;
      res_2_sum <= res_2_sum + score_2_x30;
      res_3_sum <= res_3_sum + score_3_x30;
      res_4_sum <= res_4_sum + score_4_x30;
      res_5_sum <= res_5_sum + score_5_x30;
      res_6_sum <= res_6_sum + score_6_x30;
      res_7_sum <= res_7_sum + score_7_x30;
      res_8_sum <= res_8_sum + score_8_x30;
      res_9_sum <= res_9_sum + score_9_x30;
   end
   else if(res_done_x31) begin
      res_0_sum <= res_0_sum + score_0_x31;
      res_1_sum <= res_1_sum + score_1_x31;
      res_2_sum <= res_2_sum + score_2_x31;
      res_3_sum <= res_3_sum + score_3_x31;
      res_4_sum <= res_4_sum + score_4_x31;
      res_5_sum <= res_5_sum + score_5_x31;
      res_6_sum <= res_6_sum + score_6_x31;
      res_7_sum <= res_7_sum + score_7_x31;
      res_8_sum <= res_8_sum + score_8_x31;
      res_9_sum <= res_9_sum + score_9_x31;
   end
   else if(res_done_x32) begin
      res_0_sum <= res_0_sum + score_0_x32;
      res_1_sum <= res_1_sum + score_1_x32;
      res_2_sum <= res_2_sum + score_2_x32;
      res_3_sum <= res_3_sum + score_3_x32;
      res_4_sum <= res_4_sum + score_4_x32;
      res_5_sum <= res_5_sum + score_5_x32;
      res_6_sum <= res_6_sum + score_6_x32;
      res_7_sum <= res_7_sum + score_7_x32;
      res_8_sum <= res_8_sum + score_8_x32;
      res_9_sum <= res_9_sum + score_9_x32;
   end
   else if(res_done_x33) begin
      res_0_sum <= res_0_sum + score_0_x33;
      res_1_sum <= res_1_sum + score_1_x33;
      res_2_sum <= res_2_sum + score_2_x33;
      res_3_sum <= res_3_sum + score_3_x33;
      res_4_sum <= res_4_sum + score_4_x33;
      res_5_sum <= res_5_sum + score_5_x33;
      res_6_sum <= res_6_sum + score_6_x33;
      res_7_sum <= res_7_sum + score_7_x33;
      res_8_sum <= res_8_sum + score_8_x33;
      res_9_sum <= res_9_sum + score_9_x33;
   end
   else if(res_done_x34) begin
      res_0_sum <= res_0_sum + score_0_x34;
      res_1_sum <= res_1_sum + score_1_x34;
      res_2_sum <= res_2_sum + score_2_x34;
      res_3_sum <= res_3_sum + score_3_x34;
      res_4_sum <= res_4_sum + score_4_x34;
      res_5_sum <= res_5_sum + score_5_x34;
      res_6_sum <= res_6_sum + score_6_x34;
      res_7_sum <= res_7_sum + score_7_x34;
      res_8_sum <= res_8_sum + score_8_x34;
      res_9_sum <= res_9_sum + score_9_x34;
   end
   else if(res_done_x35) begin
      res_0_sum <= res_0_sum + score_0_x35;
      res_1_sum <= res_1_sum + score_1_x35;
      res_2_sum <= res_2_sum + score_2_x35;
      res_3_sum <= res_3_sum + score_3_x35;
      res_4_sum <= res_4_sum + score_4_x35;
      res_5_sum <= res_5_sum + score_5_x35;
      res_6_sum <= res_6_sum + score_6_x35;
      res_7_sum <= res_7_sum + score_7_x35;
      res_8_sum <= res_8_sum + score_8_x35;
      res_9_sum <= res_9_sum + score_9_x35;
   end
   else if(res_done_x36) begin
      res_0_sum <= res_0_sum + score_0_x36;
      res_1_sum <= res_1_sum + score_1_x36;
      res_2_sum <= res_2_sum + score_2_x36;
      res_3_sum <= res_3_sum + score_3_x36;
      res_4_sum <= res_4_sum + score_4_x36;
      res_5_sum <= res_5_sum + score_5_x36;
      res_6_sum <= res_6_sum + score_6_x36;
      res_7_sum <= res_7_sum + score_7_x36;
      res_8_sum <= res_8_sum + score_8_x36;
      res_9_sum <= res_9_sum + score_9_x36;
   end
   else if(res_done_x37) begin
      res_0_sum <= res_0_sum + score_0_x37;
      res_1_sum <= res_1_sum + score_1_x37;
      res_2_sum <= res_2_sum + score_2_x37;
      res_3_sum <= res_3_sum + score_3_x37;
      res_4_sum <= res_4_sum + score_4_x37;
      res_5_sum <= res_5_sum + score_5_x37;
      res_6_sum <= res_6_sum + score_6_x37;
      res_7_sum <= res_7_sum + score_7_x37;
      res_8_sum <= res_8_sum + score_8_x37;
      res_9_sum <= res_9_sum + score_9_x37;
   end
   else if(res_done_x38) begin
      res_0_sum <= res_0_sum + score_0_x38;
      res_1_sum <= res_1_sum + score_1_x38;
      res_2_sum <= res_2_sum + score_2_x38;
      res_3_sum <= res_3_sum + score_3_x38;
      res_4_sum <= res_4_sum + score_4_x38;
      res_5_sum <= res_5_sum + score_5_x38;
      res_6_sum <= res_6_sum + score_6_x38;
      res_7_sum <= res_7_sum + score_7_x38;
      res_8_sum <= res_8_sum + score_8_x38;
      res_9_sum <= res_9_sum + score_9_x38;
   end
   else if(res_done_x39) begin
      res_0_sum <= res_0_sum + score_0_x39;
      res_1_sum <= res_1_sum + score_1_x39;
      res_2_sum <= res_2_sum + score_2_x39;
      res_3_sum <= res_3_sum + score_3_x39;
      res_4_sum <= res_4_sum + score_4_x39;
      res_5_sum <= res_5_sum + score_5_x39;
      res_6_sum <= res_6_sum + score_6_x39;
      res_7_sum <= res_7_sum + score_7_x39;
      res_8_sum <= res_8_sum + score_8_x39;
      res_9_sum <= res_9_sum + score_9_x39;
   end
   else if(res_done_x40) begin
      res_0_sum <= res_0_sum + score_0_x40;
      res_1_sum <= res_1_sum + score_1_x40;
      res_2_sum <= res_2_sum + score_2_x40;
      res_3_sum <= res_3_sum + score_3_x40;
      res_4_sum <= res_4_sum + score_4_x40;
      res_5_sum <= res_5_sum + score_5_x40;
      res_6_sum <= res_6_sum + score_6_x40;
      res_7_sum <= res_7_sum + score_7_x40;
      res_8_sum <= res_8_sum + score_8_x40;
      res_9_sum <= res_9_sum + score_9_x40;
   end
   else if(res_done_x41) begin
      res_0_sum <= res_0_sum + score_0_x41;
      res_1_sum <= res_1_sum + score_1_x41;
      res_2_sum <= res_2_sum + score_2_x41;
      res_3_sum <= res_3_sum + score_3_x41;
      res_4_sum <= res_4_sum + score_4_x41;
      res_5_sum <= res_5_sum + score_5_x41;
      res_6_sum <= res_6_sum + score_6_x41;
      res_7_sum <= res_7_sum + score_7_x41;
      res_8_sum <= res_8_sum + score_8_x41;
      res_9_sum <= res_9_sum + score_9_x41;
   end
   else if(res_done_x42) begin
      res_0_sum <= res_0_sum + score_0_x42;
      res_1_sum <= res_1_sum + score_1_x42;
      res_2_sum <= res_2_sum + score_2_x42;
      res_3_sum <= res_3_sum + score_3_x42;
      res_4_sum <= res_4_sum + score_4_x42;
      res_5_sum <= res_5_sum + score_5_x42;
      res_6_sum <= res_6_sum + score_6_x42;
      res_7_sum <= res_7_sum + score_7_x42;
      res_8_sum <= res_8_sum + score_8_x42;
      res_9_sum <= res_9_sum + score_9_x42;
   end
   else if(res_done_x43) begin
      res_0_sum <= res_0_sum + score_0_x43;
      res_1_sum <= res_1_sum + score_1_x43;
      res_2_sum <= res_2_sum + score_2_x43;
      res_3_sum <= res_3_sum + score_3_x43;
      res_4_sum <= res_4_sum + score_4_x43;
      res_5_sum <= res_5_sum + score_5_x43;
      res_6_sum <= res_6_sum + score_6_x43;
      res_7_sum <= res_7_sum + score_7_x43;
      res_8_sum <= res_8_sum + score_8_x43;
      res_9_sum <= res_9_sum + score_9_x43;
   end
   else if(res_done_x44) begin
      res_0_sum <= res_0_sum + score_0_x44;
      res_1_sum <= res_1_sum + score_1_x44;
      res_2_sum <= res_2_sum + score_2_x44;
      res_3_sum <= res_3_sum + score_3_x44;
      res_4_sum <= res_4_sum + score_4_x44;
      res_5_sum <= res_5_sum + score_5_x44;
      res_6_sum <= res_6_sum + score_6_x44;
      res_7_sum <= res_7_sum + score_7_x44;
      res_8_sum <= res_8_sum + score_8_x44;
      res_9_sum <= res_9_sum + score_9_x44;
   end
   else if(res_done_x45) begin
      res_0_sum <= res_0_sum + score_0_x45;
      res_1_sum <= res_1_sum + score_1_x45;
      res_2_sum <= res_2_sum + score_2_x45;
      res_3_sum <= res_3_sum + score_3_x45;
      res_4_sum <= res_4_sum + score_4_x45;
      res_5_sum <= res_5_sum + score_5_x45;
      res_6_sum <= res_6_sum + score_6_x45;
      res_7_sum <= res_7_sum + score_7_x45;
      res_8_sum <= res_8_sum + score_8_x45;
      res_9_sum <= res_9_sum + score_9_x45;
   end
   else if(res_done_x46) begin
      res_0_sum <= res_0_sum + score_0_x46;
      res_1_sum <= res_1_sum + score_1_x46;
      res_2_sum <= res_2_sum + score_2_x46;
      res_3_sum <= res_3_sum + score_3_x46;
      res_4_sum <= res_4_sum + score_4_x46;
      res_5_sum <= res_5_sum + score_5_x46;
      res_6_sum <= res_6_sum + score_6_x46;
      res_7_sum <= res_7_sum + score_7_x46;
      res_8_sum <= res_8_sum + score_8_x46;
      res_9_sum <= res_9_sum + score_9_x46;
   end
   else if(res_done_x47) begin
      res_0_sum <= res_0_sum + score_0_x47;
      res_1_sum <= res_1_sum + score_1_x47;
      res_2_sum <= res_2_sum + score_2_x47;
      res_3_sum <= res_3_sum + score_3_x47;
      res_4_sum <= res_4_sum + score_4_x47;
      res_5_sum <= res_5_sum + score_5_x47;
      res_6_sum <= res_6_sum + score_6_x47;
      res_7_sum <= res_7_sum + score_7_x47;
      res_8_sum <= res_8_sum + score_8_x47;
      res_9_sum <= res_9_sum + score_9_x47;
   end
   else if(res_done_x48) begin
      res_0_sum <= res_0_sum + score_0_x48;
      res_1_sum <= res_1_sum + score_1_x48;
      res_2_sum <= res_2_sum + score_2_x48;
      res_3_sum <= res_3_sum + score_3_x48;
      res_4_sum <= res_4_sum + score_4_x48;
      res_5_sum <= res_5_sum + score_5_x48;
      res_6_sum <= res_6_sum + score_6_x48;
      res_7_sum <= res_7_sum + score_7_x48;
      res_8_sum <= res_8_sum + score_8_x48;
      res_9_sum <= res_9_sum + score_9_x48;
   end
   else if(res_done_x49) begin
      res_0_sum <= res_0_sum + score_0_x49;
      res_1_sum <= res_1_sum + score_1_x49;
      res_2_sum <= res_2_sum + score_2_x49;
      res_3_sum <= res_3_sum + score_3_x49;
      res_4_sum <= res_4_sum + score_4_x49;
      res_5_sum <= res_5_sum + score_5_x49;
      res_6_sum <= res_6_sum + score_6_x49;
      res_7_sum <= res_7_sum + score_7_x49;
      res_8_sum <= res_8_sum + score_8_x49;
      res_9_sum <= res_9_sum + score_9_x49;
   end
   else if(res_done_x50) begin
      res_0_sum <= res_0_sum + score_0_x50;
      res_1_sum <= res_1_sum + score_1_x50;
      res_2_sum <= res_2_sum + score_2_x50;
      res_3_sum <= res_3_sum + score_3_x50;
      res_4_sum <= res_4_sum + score_4_x50;
      res_5_sum <= res_5_sum + score_5_x50;
      res_6_sum <= res_6_sum + score_6_x50;
      res_7_sum <= res_7_sum + score_7_x50;
      res_8_sum <= res_8_sum + score_8_x50;
      res_9_sum <= res_9_sum + score_9_x50;
   end
   else if(res_done_x51) begin
      res_0_sum <= res_0_sum + score_0_x51;
      res_1_sum <= res_1_sum + score_1_x51;
      res_2_sum <= res_2_sum + score_2_x51;
      res_3_sum <= res_3_sum + score_3_x51;
      res_4_sum <= res_4_sum + score_4_x51;
      res_5_sum <= res_5_sum + score_5_x51;
      res_6_sum <= res_6_sum + score_6_x51;
      res_7_sum <= res_7_sum + score_7_x51;
      res_8_sum <= res_8_sum + score_8_x51;
      res_9_sum <= res_9_sum + score_9_x51;
   end
   else if(res_done_x52) begin
      res_0_sum <= res_0_sum + score_0_x52;
      res_1_sum <= res_1_sum + score_1_x52;
      res_2_sum <= res_2_sum + score_2_x52;
      res_3_sum <= res_3_sum + score_3_x52;
      res_4_sum <= res_4_sum + score_4_x52;
      res_5_sum <= res_5_sum + score_5_x52;
      res_6_sum <= res_6_sum + score_6_x52;
      res_7_sum <= res_7_sum + score_7_x52;
      res_8_sum <= res_8_sum + score_8_x52;
      res_9_sum <= res_9_sum + score_9_x52;
   end
   else if(res_done_x53) begin
      res_0_sum <= res_0_sum + score_0_x53;
      res_1_sum <= res_1_sum + score_1_x53;
      res_2_sum <= res_2_sum + score_2_x53;
      res_3_sum <= res_3_sum + score_3_x53;
      res_4_sum <= res_4_sum + score_4_x53;
      res_5_sum <= res_5_sum + score_5_x53;
      res_6_sum <= res_6_sum + score_6_x53;
      res_7_sum <= res_7_sum + score_7_x53;
      res_8_sum <= res_8_sum + score_8_x53;
      res_9_sum <= res_9_sum + score_9_x53;
   end
   else if(res_done_x54) begin
      res_0_sum <= res_0_sum + score_0_x54;
      res_1_sum <= res_1_sum + score_1_x54;
      res_2_sum <= res_2_sum + score_2_x54;
      res_3_sum <= res_3_sum + score_3_x54;
      res_4_sum <= res_4_sum + score_4_x54;
      res_5_sum <= res_5_sum + score_5_x54;
      res_6_sum <= res_6_sum + score_6_x54;
      res_7_sum <= res_7_sum + score_7_x54;
      res_8_sum <= res_8_sum + score_8_x54;
      res_9_sum <= res_9_sum + score_9_x54;
   end
   else if(res_done_x55) begin
      res_0_sum <= res_0_sum + score_0_x55;
      res_1_sum <= res_1_sum + score_1_x55;
      res_2_sum <= res_2_sum + score_2_x55;
      res_3_sum <= res_3_sum + score_3_x55;
      res_4_sum <= res_4_sum + score_4_x55;
      res_5_sum <= res_5_sum + score_5_x55;
      res_6_sum <= res_6_sum + score_6_x55;
      res_7_sum <= res_7_sum + score_7_x55;
      res_8_sum <= res_8_sum + score_8_x55;
      res_9_sum <= res_9_sum + score_9_x55;
   end
   else if(res_done_x56) begin
      res_0_sum <= res_0_sum + score_0_x56;
      res_1_sum <= res_1_sum + score_1_x56;
      res_2_sum <= res_2_sum + score_2_x56;
      res_3_sum <= res_3_sum + score_3_x56;
      res_4_sum <= res_4_sum + score_4_x56;
      res_5_sum <= res_5_sum + score_5_x56;
      res_6_sum <= res_6_sum + score_6_x56;
      res_7_sum <= res_7_sum + score_7_x56;
      res_8_sum <= res_8_sum + score_8_x56;
      res_9_sum <= res_9_sum + score_9_x56;
   end
   else if(res_done_x57) begin
      res_0_sum <= res_0_sum + score_0_x57;
      res_1_sum <= res_1_sum + score_1_x57;
      res_2_sum <= res_2_sum + score_2_x57;
      res_3_sum <= res_3_sum + score_3_x57;
      res_4_sum <= res_4_sum + score_4_x57;
      res_5_sum <= res_5_sum + score_5_x57;
      res_6_sum <= res_6_sum + score_6_x57;
      res_7_sum <= res_7_sum + score_7_x57;
      res_8_sum <= res_8_sum + score_8_x57;
      res_9_sum <= res_9_sum + score_9_x57;
   end
   else if(res_done_x58) begin
      res_0_sum <= res_0_sum + score_0_x58;
      res_1_sum <= res_1_sum + score_1_x58;
      res_2_sum <= res_2_sum + score_2_x58;
      res_3_sum <= res_3_sum + score_3_x58;
      res_4_sum <= res_4_sum + score_4_x58;
      res_5_sum <= res_5_sum + score_5_x58;
      res_6_sum <= res_6_sum + score_6_x58;
      res_7_sum <= res_7_sum + score_7_x58;
      res_8_sum <= res_8_sum + score_8_x58;
      res_9_sum <= res_9_sum + score_9_x58;
   end
   else if(res_done_x59) begin
      res_0_sum <= res_0_sum + score_0_x59;
      res_1_sum <= res_1_sum + score_1_x59;
      res_2_sum <= res_2_sum + score_2_x59;
      res_3_sum <= res_3_sum + score_3_x59;
      res_4_sum <= res_4_sum + score_4_x59;
      res_5_sum <= res_5_sum + score_5_x59;
      res_6_sum <= res_6_sum + score_6_x59;
      res_7_sum <= res_7_sum + score_7_x59;
      res_8_sum <= res_8_sum + score_8_x59;
      res_9_sum <= res_9_sum + score_9_x59;
   end
   else if(res_done_x60) begin
      res_0_sum <= res_0_sum + score_0_x60;
      res_1_sum <= res_1_sum + score_1_x60;
      res_2_sum <= res_2_sum + score_2_x60;
      res_3_sum <= res_3_sum + score_3_x60;
      res_4_sum <= res_4_sum + score_4_x60;
      res_5_sum <= res_5_sum + score_5_x60;
      res_6_sum <= res_6_sum + score_6_x60;
      res_7_sum <= res_7_sum + score_7_x60;
      res_8_sum <= res_8_sum + score_8_x60;
      res_9_sum <= res_9_sum + score_9_x60;
   end
   else if(res_done_x61) begin
      res_0_sum <= res_0_sum + score_0_x61;
      res_1_sum <= res_1_sum + score_1_x61;
      res_2_sum <= res_2_sum + score_2_x61;
      res_3_sum <= res_3_sum + score_3_x61;
      res_4_sum <= res_4_sum + score_4_x61;
      res_5_sum <= res_5_sum + score_5_x61;
      res_6_sum <= res_6_sum + score_6_x61;
      res_7_sum <= res_7_sum + score_7_x61;
      res_8_sum <= res_8_sum + score_8_x61;
      res_9_sum <= res_9_sum + score_9_x61;
   end
   else if(res_done_x62) begin
      res_0_sum <= res_0_sum + score_0_x62;
      res_1_sum <= res_1_sum + score_1_x62;
      res_2_sum <= res_2_sum + score_2_x62;
      res_3_sum <= res_3_sum + score_3_x62;
      res_4_sum <= res_4_sum + score_4_x62;
      res_5_sum <= res_5_sum + score_5_x62;
      res_6_sum <= res_6_sum + score_6_x62;
      res_7_sum <= res_7_sum + score_7_x62;
      res_8_sum <= res_8_sum + score_8_x62;
      res_9_sum <= res_9_sum + score_9_x62;
   end
   else if(res_done_x63) begin
      res_0_sum <= res_0_sum + score_0_x63;
      res_1_sum <= res_1_sum + score_1_x63;
      res_2_sum <= res_2_sum + score_2_x63;
      res_3_sum <= res_3_sum + score_3_x63;
      res_4_sum <= res_4_sum + score_4_x63;
      res_5_sum <= res_5_sum + score_5_x63;
      res_6_sum <= res_6_sum + score_6_x63;
      res_7_sum <= res_7_sum + score_7_x63;
      res_8_sum <= res_8_sum + score_8_x63;
      res_9_sum <= res_9_sum + score_9_x63;
   end
   else if(res_done_x64) begin
      res_0_sum <= res_0_sum + score_0_x64;
      res_1_sum <= res_1_sum + score_1_x64;
      res_2_sum <= res_2_sum + score_2_x64;
      res_3_sum <= res_3_sum + score_3_x64;
      res_4_sum <= res_4_sum + score_4_x64;
      res_5_sum <= res_5_sum + score_5_x64;
      res_6_sum <= res_6_sum + score_6_x64;
      res_7_sum <= res_7_sum + score_7_x64;
      res_8_sum <= res_8_sum + score_8_x64;
      res_9_sum <= res_9_sum + score_9_x64;
   end
   else if(res_done_x65) begin
      res_0_sum <= res_0_sum + score_0_x65;
      res_1_sum <= res_1_sum + score_1_x65;
      res_2_sum <= res_2_sum + score_2_x65;
      res_3_sum <= res_3_sum + score_3_x65;
      res_4_sum <= res_4_sum + score_4_x65;
      res_5_sum <= res_5_sum + score_5_x65;
      res_6_sum <= res_6_sum + score_6_x65;
      res_7_sum <= res_7_sum + score_7_x65;
      res_8_sum <= res_8_sum + score_8_x65;
      res_9_sum <= res_9_sum + score_9_x65;
   end
   else if(res_done_x66) begin
      res_0_sum <= res_0_sum + score_0_x66;
      res_1_sum <= res_1_sum + score_1_x66;
      res_2_sum <= res_2_sum + score_2_x66;
      res_3_sum <= res_3_sum + score_3_x66;
      res_4_sum <= res_4_sum + score_4_x66;
      res_5_sum <= res_5_sum + score_5_x66;
      res_6_sum <= res_6_sum + score_6_x66;
      res_7_sum <= res_7_sum + score_7_x66;
      res_8_sum <= res_8_sum + score_8_x66;
      res_9_sum <= res_9_sum + score_9_x66;
   end
   else if(res_done_x67) begin
      res_0_sum <= res_0_sum + score_0_x67;
      res_1_sum <= res_1_sum + score_1_x67;
      res_2_sum <= res_2_sum + score_2_x67;
      res_3_sum <= res_3_sum + score_3_x67;
      res_4_sum <= res_4_sum + score_4_x67;
      res_5_sum <= res_5_sum + score_5_x67;
      res_6_sum <= res_6_sum + score_6_x67;
      res_7_sum <= res_7_sum + score_7_x67;
      res_8_sum <= res_8_sum + score_8_x67;
      res_9_sum <= res_9_sum + score_9_x67;
   end
   else if(res_done_x68) begin
      res_0_sum <= res_0_sum + score_0_x68;
      res_1_sum <= res_1_sum + score_1_x68;
      res_2_sum <= res_2_sum + score_2_x68;
      res_3_sum <= res_3_sum + score_3_x68;
      res_4_sum <= res_4_sum + score_4_x68;
      res_5_sum <= res_5_sum + score_5_x68;
      res_6_sum <= res_6_sum + score_6_x68;
      res_7_sum <= res_7_sum + score_7_x68;
      res_8_sum <= res_8_sum + score_8_x68;
      res_9_sum <= res_9_sum + score_9_x68;
   end
   else if(res_done_x69) begin
      res_0_sum <= res_0_sum + score_0_x69;
      res_1_sum <= res_1_sum + score_1_x69;
      res_2_sum <= res_2_sum + score_2_x69;
      res_3_sum <= res_3_sum + score_3_x69;
      res_4_sum <= res_4_sum + score_4_x69;
      res_5_sum <= res_5_sum + score_5_x69;
      res_6_sum <= res_6_sum + score_6_x69;
      res_7_sum <= res_7_sum + score_7_x69;
      res_8_sum <= res_8_sum + score_8_x69;
      res_9_sum <= res_9_sum + score_9_x69;
   end
   else if(res_done_x70) begin
      res_0_sum <= res_0_sum + score_0_x70;
      res_1_sum <= res_1_sum + score_1_x70;
      res_2_sum <= res_2_sum + score_2_x70;
      res_3_sum <= res_3_sum + score_3_x70;
      res_4_sum <= res_4_sum + score_4_x70;
      res_5_sum <= res_5_sum + score_5_x70;
      res_6_sum <= res_6_sum + score_6_x70;
      res_7_sum <= res_7_sum + score_7_x70;
      res_8_sum <= res_8_sum + score_8_x70;
      res_9_sum <= res_9_sum + score_9_x70;
   end
   else if(res_done_x71) begin
      res_0_sum <= res_0_sum + score_0_x71;
      res_1_sum <= res_1_sum + score_1_x71;
      res_2_sum <= res_2_sum + score_2_x71;
      res_3_sum <= res_3_sum + score_3_x71;
      res_4_sum <= res_4_sum + score_4_x71;
      res_5_sum <= res_5_sum + score_5_x71;
      res_6_sum <= res_6_sum + score_6_x71;
      res_7_sum <= res_7_sum + score_7_x71;
      res_8_sum <= res_8_sum + score_8_x71;
      res_9_sum <= res_9_sum + score_9_x71;
   end
   else if(res_done_x72) begin
      res_0_sum <= res_0_sum + score_0_x72;
      res_1_sum <= res_1_sum + score_1_x72;
      res_2_sum <= res_2_sum + score_2_x72;
      res_3_sum <= res_3_sum + score_3_x72;
      res_4_sum <= res_4_sum + score_4_x72;
      res_5_sum <= res_5_sum + score_5_x72;
      res_6_sum <= res_6_sum + score_6_x72;
      res_7_sum <= res_7_sum + score_7_x72;
      res_8_sum <= res_8_sum + score_8_x72;
      res_9_sum <= res_9_sum + score_9_x72;
   end
   else if(res_done_x73) begin
      res_0_sum <= res_0_sum + score_0_x73;
      res_1_sum <= res_1_sum + score_1_x73;
      res_2_sum <= res_2_sum + score_2_x73;
      res_3_sum <= res_3_sum + score_3_x73;
      res_4_sum <= res_4_sum + score_4_x73;
      res_5_sum <= res_5_sum + score_5_x73;
      res_6_sum <= res_6_sum + score_6_x73;
      res_7_sum <= res_7_sum + score_7_x73;
      res_8_sum <= res_8_sum + score_8_x73;
      res_9_sum <= res_9_sum + score_9_x73;
   end
   else if(res_done_x74) begin
      res_0_sum <= res_0_sum + score_0_x74;
      res_1_sum <= res_1_sum + score_1_x74;
      res_2_sum <= res_2_sum + score_2_x74;
      res_3_sum <= res_3_sum + score_3_x74;
      res_4_sum <= res_4_sum + score_4_x74;
      res_5_sum <= res_5_sum + score_5_x74;
      res_6_sum <= res_6_sum + score_6_x74;
      res_7_sum <= res_7_sum + score_7_x74;
      res_8_sum <= res_8_sum + score_8_x74;
      res_9_sum <= res_9_sum + score_9_x74;
   end
   else if(res_done_x75) begin
      res_0_sum <= res_0_sum + score_0_x75;
      res_1_sum <= res_1_sum + score_1_x75;
      res_2_sum <= res_2_sum + score_2_x75;
      res_3_sum <= res_3_sum + score_3_x75;
      res_4_sum <= res_4_sum + score_4_x75;
      res_5_sum <= res_5_sum + score_5_x75;
      res_6_sum <= res_6_sum + score_6_x75;
      res_7_sum <= res_7_sum + score_7_x75;
      res_8_sum <= res_8_sum + score_8_x75;
      res_9_sum <= res_9_sum + score_9_x75;
   end
   else if(res_done_x76) begin
      res_0_sum <= res_0_sum + score_0_x76;
      res_1_sum <= res_1_sum + score_1_x76;
      res_2_sum <= res_2_sum + score_2_x76;
      res_3_sum <= res_3_sum + score_3_x76;
      res_4_sum <= res_4_sum + score_4_x76;
      res_5_sum <= res_5_sum + score_5_x76;
      res_6_sum <= res_6_sum + score_6_x76;
      res_7_sum <= res_7_sum + score_7_x76;
      res_8_sum <= res_8_sum + score_8_x76;
      res_9_sum <= res_9_sum + score_9_x76;
   end
   else if(res_done_x77) begin
      res_0_sum <= res_0_sum + score_0_x77;
      res_1_sum <= res_1_sum + score_1_x77;
      res_2_sum <= res_2_sum + score_2_x77;
      res_3_sum <= res_3_sum + score_3_x77;
      res_4_sum <= res_4_sum + score_4_x77;
      res_5_sum <= res_5_sum + score_5_x77;
      res_6_sum <= res_6_sum + score_6_x77;
      res_7_sum <= res_7_sum + score_7_x77;
      res_8_sum <= res_8_sum + score_8_x77;
      res_9_sum <= res_9_sum + score_9_x77;
   end
   else if(res_done_x78) begin
      res_0_sum <= res_0_sum + score_0_x78;
      res_1_sum <= res_1_sum + score_1_x78;
      res_2_sum <= res_2_sum + score_2_x78;
      res_3_sum <= res_3_sum + score_3_x78;
      res_4_sum <= res_4_sum + score_4_x78;
      res_5_sum <= res_5_sum + score_5_x78;
      res_6_sum <= res_6_sum + score_6_x78;
      res_7_sum <= res_7_sum + score_7_x78;
      res_8_sum <= res_8_sum + score_8_x78;
      res_9_sum <= res_9_sum + score_9_x78;
   end
   else if(res_done_x79) begin
      res_0_sum <= res_0_sum + score_0_x79;
      res_1_sum <= res_1_sum + score_1_x79;
      res_2_sum <= res_2_sum + score_2_x79;
      res_3_sum <= res_3_sum + score_3_x79;
      res_4_sum <= res_4_sum + score_4_x79;
      res_5_sum <= res_5_sum + score_5_x79;
      res_6_sum <= res_6_sum + score_6_x79;
      res_7_sum <= res_7_sum + score_7_x79;
      res_8_sum <= res_8_sum + score_8_x79;
      res_9_sum <= res_9_sum + score_9_x79;
   end
   else if(res_done_x80) begin
      res_0_sum <= res_0_sum + score_0_x80;
      res_1_sum <= res_1_sum + score_1_x80;
      res_2_sum <= res_2_sum + score_2_x80;
      res_3_sum <= res_3_sum + score_3_x80;
      res_4_sum <= res_4_sum + score_4_x80;
      res_5_sum <= res_5_sum + score_5_x80;
      res_6_sum <= res_6_sum + score_6_x80;
      res_7_sum <= res_7_sum + score_7_x80;
      res_8_sum <= res_8_sum + score_8_x80;
      res_9_sum <= res_9_sum + score_9_x80;
   end
   else if(res_done_x81) begin
      res_0_sum <= res_0_sum + score_0_x81;
      res_1_sum <= res_1_sum + score_1_x81;
      res_2_sum <= res_2_sum + score_2_x81;
      res_3_sum <= res_3_sum + score_3_x81;
      res_4_sum <= res_4_sum + score_4_x81;
      res_5_sum <= res_5_sum + score_5_x81;
      res_6_sum <= res_6_sum + score_6_x81;
      res_7_sum <= res_7_sum + score_7_x81;
      res_8_sum <= res_8_sum + score_8_x81;
      res_9_sum <= res_9_sum + score_9_x81;
   end
   else if(res_done_x82) begin
      res_0_sum <= res_0_sum + score_0_x82;
      res_1_sum <= res_1_sum + score_1_x82;
      res_2_sum <= res_2_sum + score_2_x82;
      res_3_sum <= res_3_sum + score_3_x82;
      res_4_sum <= res_4_sum + score_4_x82;
      res_5_sum <= res_5_sum + score_5_x82;
      res_6_sum <= res_6_sum + score_6_x82;
      res_7_sum <= res_7_sum + score_7_x82;
      res_8_sum <= res_8_sum + score_8_x82;
      res_9_sum <= res_9_sum + score_9_x82;
   end
   else if(res_done_x83) begin
      res_0_sum <= res_0_sum + score_0_x83;
      res_1_sum <= res_1_sum + score_1_x83;
      res_2_sum <= res_2_sum + score_2_x83;
      res_3_sum <= res_3_sum + score_3_x83;
      res_4_sum <= res_4_sum + score_4_x83;
      res_5_sum <= res_5_sum + score_5_x83;
      res_6_sum <= res_6_sum + score_6_x83;
      res_7_sum <= res_7_sum + score_7_x83;
      res_8_sum <= res_8_sum + score_8_x83;
      res_9_sum <= res_9_sum + score_9_x83;
   end
   else if(res_done_x84) begin
      res_0_sum <= res_0_sum + score_0_x84;
      res_1_sum <= res_1_sum + score_1_x84;
      res_2_sum <= res_2_sum + score_2_x84;
      res_3_sum <= res_3_sum + score_3_x84;
      res_4_sum <= res_4_sum + score_4_x84;
      res_5_sum <= res_5_sum + score_5_x84;
      res_6_sum <= res_6_sum + score_6_x84;
      res_7_sum <= res_7_sum + score_7_x84;
      res_8_sum <= res_8_sum + score_8_x84;
      res_9_sum <= res_9_sum + score_9_x84;
   end
   else if(res_done_x85) begin
      res_0_sum <= res_0_sum + score_0_x85;
      res_1_sum <= res_1_sum + score_1_x85;
      res_2_sum <= res_2_sum + score_2_x85;
      res_3_sum <= res_3_sum + score_3_x85;
      res_4_sum <= res_4_sum + score_4_x85;
      res_5_sum <= res_5_sum + score_5_x85;
      res_6_sum <= res_6_sum + score_6_x85;
      res_7_sum <= res_7_sum + score_7_x85;
      res_8_sum <= res_8_sum + score_8_x85;
      res_9_sum <= res_9_sum + score_9_x85;
   end
   else if(res_done_x86) begin
      res_0_sum <= res_0_sum + score_0_x86;
      res_1_sum <= res_1_sum + score_1_x86;
      res_2_sum <= res_2_sum + score_2_x86;
      res_3_sum <= res_3_sum + score_3_x86;
      res_4_sum <= res_4_sum + score_4_x86;
      res_5_sum <= res_5_sum + score_5_x86;
      res_6_sum <= res_6_sum + score_6_x86;
      res_7_sum <= res_7_sum + score_7_x86;
      res_8_sum <= res_8_sum + score_8_x86;
      res_9_sum <= res_9_sum + score_9_x86;
   end
   else if(res_done_x87) begin
      res_0_sum <= res_0_sum + score_0_x87;
      res_1_sum <= res_1_sum + score_1_x87;
      res_2_sum <= res_2_sum + score_2_x87;
      res_3_sum <= res_3_sum + score_3_x87;
      res_4_sum <= res_4_sum + score_4_x87;
      res_5_sum <= res_5_sum + score_5_x87;
      res_6_sum <= res_6_sum + score_6_x87;
      res_7_sum <= res_7_sum + score_7_x87;
      res_8_sum <= res_8_sum + score_8_x87;
      res_9_sum <= res_9_sum + score_9_x87;
   end
   else if(res_done_x88) begin
      res_0_sum <= res_0_sum + score_0_x88;
      res_1_sum <= res_1_sum + score_1_x88;
      res_2_sum <= res_2_sum + score_2_x88;
      res_3_sum <= res_3_sum + score_3_x88;
      res_4_sum <= res_4_sum + score_4_x88;
      res_5_sum <= res_5_sum + score_5_x88;
      res_6_sum <= res_6_sum + score_6_x88;
      res_7_sum <= res_7_sum + score_7_x88;
      res_8_sum <= res_8_sum + score_8_x88;
      res_9_sum <= res_9_sum + score_9_x88;
   end
   else if(res_done_x89) begin
      res_0_sum <= res_0_sum + score_0_x89;
      res_1_sum <= res_1_sum + score_1_x89;
      res_2_sum <= res_2_sum + score_2_x89;
      res_3_sum <= res_3_sum + score_3_x89;
      res_4_sum <= res_4_sum + score_4_x89;
      res_5_sum <= res_5_sum + score_5_x89;
      res_6_sum <= res_6_sum + score_6_x89;
      res_7_sum <= res_7_sum + score_7_x89;
      res_8_sum <= res_8_sum + score_8_x89;
      res_9_sum <= res_9_sum + score_9_x89;
   end
   else if(res_done_x90) begin
      res_0_sum <= res_0_sum + score_0_x90;
      res_1_sum <= res_1_sum + score_1_x90;
      res_2_sum <= res_2_sum + score_2_x90;
      res_3_sum <= res_3_sum + score_3_x90;
      res_4_sum <= res_4_sum + score_4_x90;
      res_5_sum <= res_5_sum + score_5_x90;
      res_6_sum <= res_6_sum + score_6_x90;
      res_7_sum <= res_7_sum + score_7_x90;
      res_8_sum <= res_8_sum + score_8_x90;
      res_9_sum <= res_9_sum + score_9_x90;
   end
   else if(res_done_x91) begin
      res_0_sum <= res_0_sum + score_0_x91;
      res_1_sum <= res_1_sum + score_1_x91;
      res_2_sum <= res_2_sum + score_2_x91;
      res_3_sum <= res_3_sum + score_3_x91;
      res_4_sum <= res_4_sum + score_4_x91;
      res_5_sum <= res_5_sum + score_5_x91;
      res_6_sum <= res_6_sum + score_6_x91;
      res_7_sum <= res_7_sum + score_7_x91;
      res_8_sum <= res_8_sum + score_8_x91;
      res_9_sum <= res_9_sum + score_9_x91;
   end
   else if(res_done_x92) begin
      res_0_sum <= res_0_sum + score_0_x92;
      res_1_sum <= res_1_sum + score_1_x92;
      res_2_sum <= res_2_sum + score_2_x92;
      res_3_sum <= res_3_sum + score_3_x92;
      res_4_sum <= res_4_sum + score_4_x92;
      res_5_sum <= res_5_sum + score_5_x92;
      res_6_sum <= res_6_sum + score_6_x92;
      res_7_sum <= res_7_sum + score_7_x92;
      res_8_sum <= res_8_sum + score_8_x92;
      res_9_sum <= res_9_sum + score_9_x92;
   end
   else if(res_done_x93) begin
      res_0_sum <= res_0_sum + score_0_x93;
      res_1_sum <= res_1_sum + score_1_x93;
      res_2_sum <= res_2_sum + score_2_x93;
      res_3_sum <= res_3_sum + score_3_x93;
      res_4_sum <= res_4_sum + score_4_x93;
      res_5_sum <= res_5_sum + score_5_x93;
      res_6_sum <= res_6_sum + score_6_x93;
      res_7_sum <= res_7_sum + score_7_x93;
      res_8_sum <= res_8_sum + score_8_x93;
      res_9_sum <= res_9_sum + score_9_x93;
   end
   else if(res_done_x94) begin
      res_0_sum <= res_0_sum + score_0_x94;
      res_1_sum <= res_1_sum + score_1_x94;
      res_2_sum <= res_2_sum + score_2_x94;
      res_3_sum <= res_3_sum + score_3_x94;
      res_4_sum <= res_4_sum + score_4_x94;
      res_5_sum <= res_5_sum + score_5_x94;
      res_6_sum <= res_6_sum + score_6_x94;
      res_7_sum <= res_7_sum + score_7_x94;
      res_8_sum <= res_8_sum + score_8_x94;
      res_9_sum <= res_9_sum + score_9_x94;
   end
   else if(res_done_x95) begin
      res_0_sum <= res_0_sum + score_0_x95;
      res_1_sum <= res_1_sum + score_1_x95;
      res_2_sum <= res_2_sum + score_2_x95;
      res_3_sum <= res_3_sum + score_3_x95;
      res_4_sum <= res_4_sum + score_4_x95;
      res_5_sum <= res_5_sum + score_5_x95;
      res_6_sum <= res_6_sum + score_6_x95;
      res_7_sum <= res_7_sum + score_7_x95;
      res_8_sum <= res_8_sum + score_8_x95;
      res_9_sum <= res_9_sum + score_9_x95;
   end
   else if(res_done_x96) begin
      res_0_sum <= res_0_sum + score_0_x96;
      res_1_sum <= res_1_sum + score_1_x96;
      res_2_sum <= res_2_sum + score_2_x96;
      res_3_sum <= res_3_sum + score_3_x96;
      res_4_sum <= res_4_sum + score_4_x96;
      res_5_sum <= res_5_sum + score_5_x96;
      res_6_sum <= res_6_sum + score_6_x96;
      res_7_sum <= res_7_sum + score_7_x96;
      res_8_sum <= res_8_sum + score_8_x96;
      res_9_sum <= res_9_sum + score_9_x96;
   end
   else if(res_done_x97) begin
      res_0_sum <= res_0_sum + score_0_x97;
      res_1_sum <= res_1_sum + score_1_x97;
      res_2_sum <= res_2_sum + score_2_x97;
      res_3_sum <= res_3_sum + score_3_x97;
      res_4_sum <= res_4_sum + score_4_x97;
      res_5_sum <= res_5_sum + score_5_x97;
      res_6_sum <= res_6_sum + score_6_x97;
      res_7_sum <= res_7_sum + score_7_x97;
      res_8_sum <= res_8_sum + score_8_x97;
      res_9_sum <= res_9_sum + score_9_x97;
   end
   else if(res_done_x98) begin
      res_0_sum <= res_0_sum + score_0_x98;
      res_1_sum <= res_1_sum + score_1_x98;
      res_2_sum <= res_2_sum + score_2_x98;
      res_3_sum <= res_3_sum + score_3_x98;
      res_4_sum <= res_4_sum + score_4_x98;
      res_5_sum <= res_5_sum + score_5_x98;
      res_6_sum <= res_6_sum + score_6_x98;
      res_7_sum <= res_7_sum + score_7_x98;
      res_8_sum <= res_8_sum + score_8_x98;
      res_9_sum <= res_9_sum + score_9_x98;
   end
   else if(res_done_x99) begin
      res_0_sum <= res_0_sum + score_0_x99;
      res_1_sum <= res_1_sum + score_1_x99;
      res_2_sum <= res_2_sum + score_2_x99;
      res_3_sum <= res_3_sum + score_3_x99;
      res_4_sum <= res_4_sum + score_4_x99;
      res_5_sum <= res_5_sum + score_5_x99;
      res_6_sum <= res_6_sum + score_6_x99;
      res_7_sum <= res_7_sum + score_7_x99;
      res_8_sum <= res_8_sum + score_8_x99;
      res_9_sum <= res_9_sum + score_9_x99;
   end
   else if(res_done_x100) begin
      res_0_sum <= res_0_sum + score_0_x100;
      res_1_sum <= res_1_sum + score_1_x100;
      res_2_sum <= res_2_sum + score_2_x100;
      res_3_sum <= res_3_sum + score_3_x100;
      res_4_sum <= res_4_sum + score_4_x100;
      res_5_sum <= res_5_sum + score_5_x100;
      res_6_sum <= res_6_sum + score_6_x100;
      res_7_sum <= res_7_sum + score_7_x100;
      res_8_sum <= res_8_sum + score_8_x100;
      res_9_sum <= res_9_sum + score_9_x100;
   end
   else if(res_done_x101) begin
      res_0_sum <= res_0_sum + score_0_x101;
      res_1_sum <= res_1_sum + score_1_x101;
      res_2_sum <= res_2_sum + score_2_x101;
      res_3_sum <= res_3_sum + score_3_x101;
      res_4_sum <= res_4_sum + score_4_x101;
      res_5_sum <= res_5_sum + score_5_x101;
      res_6_sum <= res_6_sum + score_6_x101;
      res_7_sum <= res_7_sum + score_7_x101;
      res_8_sum <= res_8_sum + score_8_x101;
      res_9_sum <= res_9_sum + score_9_x101;
   end
   else if(res_done_x102) begin
      res_0_sum <= res_0_sum + score_0_x102;
      res_1_sum <= res_1_sum + score_1_x102;
      res_2_sum <= res_2_sum + score_2_x102;
      res_3_sum <= res_3_sum + score_3_x102;
      res_4_sum <= res_4_sum + score_4_x102;
      res_5_sum <= res_5_sum + score_5_x102;
      res_6_sum <= res_6_sum + score_6_x102;
      res_7_sum <= res_7_sum + score_7_x102;
      res_8_sum <= res_8_sum + score_8_x102;
      res_9_sum <= res_9_sum + score_9_x102;
   end
   else if(res_done_x103) begin
      res_0_sum <= res_0_sum + score_0_x103;
      res_1_sum <= res_1_sum + score_1_x103;
      res_2_sum <= res_2_sum + score_2_x103;
      res_3_sum <= res_3_sum + score_3_x103;
      res_4_sum <= res_4_sum + score_4_x103;
      res_5_sum <= res_5_sum + score_5_x103;
      res_6_sum <= res_6_sum + score_6_x103;
      res_7_sum <= res_7_sum + score_7_x103;
      res_8_sum <= res_8_sum + score_8_x103;
      res_9_sum <= res_9_sum + score_9_x103;
   end
   else if(res_done_x104) begin
      res_0_sum <= res_0_sum + score_0_x104;
      res_1_sum <= res_1_sum + score_1_x104;
      res_2_sum <= res_2_sum + score_2_x104;
      res_3_sum <= res_3_sum + score_3_x104;
      res_4_sum <= res_4_sum + score_4_x104;
      res_5_sum <= res_5_sum + score_5_x104;
      res_6_sum <= res_6_sum + score_6_x104;
      res_7_sum <= res_7_sum + score_7_x104;
      res_8_sum <= res_8_sum + score_8_x104;
      res_9_sum <= res_9_sum + score_9_x104;
   end
   else if(res_done_x105) begin
      res_0_sum <= res_0_sum + score_0_x105;
      res_1_sum <= res_1_sum + score_1_x105;
      res_2_sum <= res_2_sum + score_2_x105;
      res_3_sum <= res_3_sum + score_3_x105;
      res_4_sum <= res_4_sum + score_4_x105;
      res_5_sum <= res_5_sum + score_5_x105;
      res_6_sum <= res_6_sum + score_6_x105;
      res_7_sum <= res_7_sum + score_7_x105;
      res_8_sum <= res_8_sum + score_8_x105;
      res_9_sum <= res_9_sum + score_9_x105;
   end
   else if(res_done_x106) begin
      res_0_sum <= res_0_sum + score_0_x106;
      res_1_sum <= res_1_sum + score_1_x106;
      res_2_sum <= res_2_sum + score_2_x106;
      res_3_sum <= res_3_sum + score_3_x106;
      res_4_sum <= res_4_sum + score_4_x106;
      res_5_sum <= res_5_sum + score_5_x106;
      res_6_sum <= res_6_sum + score_6_x106;
      res_7_sum <= res_7_sum + score_7_x106;
      res_8_sum <= res_8_sum + score_8_x106;
      res_9_sum <= res_9_sum + score_9_x106;
   end
   else if(res_done_x107) begin
      res_0_sum <= res_0_sum + score_0_x107;
      res_1_sum <= res_1_sum + score_1_x107;
      res_2_sum <= res_2_sum + score_2_x107;
      res_3_sum <= res_3_sum + score_3_x107;
      res_4_sum <= res_4_sum + score_4_x107;
      res_5_sum <= res_5_sum + score_5_x107;
      res_6_sum <= res_6_sum + score_6_x107;
      res_7_sum <= res_7_sum + score_7_x107;
      res_8_sum <= res_8_sum + score_8_x107;
      res_9_sum <= res_9_sum + score_9_x107;
   end
   else if(res_done_x108) begin
      res_0_sum <= res_0_sum + score_0_x108;
      res_1_sum <= res_1_sum + score_1_x108;
      res_2_sum <= res_2_sum + score_2_x108;
      res_3_sum <= res_3_sum + score_3_x108;
      res_4_sum <= res_4_sum + score_4_x108;
      res_5_sum <= res_5_sum + score_5_x108;
      res_6_sum <= res_6_sum + score_6_x108;
      res_7_sum <= res_7_sum + score_7_x108;
      res_8_sum <= res_8_sum + score_8_x108;
      res_9_sum <= res_9_sum + score_9_x108;
   end
   else if(res_done_x109) begin
      res_0_sum <= res_0_sum + score_0_x109;
      res_1_sum <= res_1_sum + score_1_x109;
      res_2_sum <= res_2_sum + score_2_x109;
      res_3_sum <= res_3_sum + score_3_x109;
      res_4_sum <= res_4_sum + score_4_x109;
      res_5_sum <= res_5_sum + score_5_x109;
      res_6_sum <= res_6_sum + score_6_x109;
      res_7_sum <= res_7_sum + score_7_x109;
      res_8_sum <= res_8_sum + score_8_x109;
      res_9_sum <= res_9_sum + score_9_x109;
   end
   else if(res_done_x110) begin
      res_0_sum <= res_0_sum + score_0_x110;
      res_1_sum <= res_1_sum + score_1_x110;
      res_2_sum <= res_2_sum + score_2_x110;
      res_3_sum <= res_3_sum + score_3_x110;
      res_4_sum <= res_4_sum + score_4_x110;
      res_5_sum <= res_5_sum + score_5_x110;
      res_6_sum <= res_6_sum + score_6_x110;
      res_7_sum <= res_7_sum + score_7_x110;
      res_8_sum <= res_8_sum + score_8_x110;
      res_9_sum <= res_9_sum + score_9_x110;
   end
   else if(res_done_x111) begin
      res_0_sum <= res_0_sum + score_0_x111;
      res_1_sum <= res_1_sum + score_1_x111;
      res_2_sum <= res_2_sum + score_2_x111;
      res_3_sum <= res_3_sum + score_3_x111;
      res_4_sum <= res_4_sum + score_4_x111;
      res_5_sum <= res_5_sum + score_5_x111;
      res_6_sum <= res_6_sum + score_6_x111;
      res_7_sum <= res_7_sum + score_7_x111;
      res_8_sum <= res_8_sum + score_8_x111;
      res_9_sum <= res_9_sum + score_9_x111;
   end
   else if(res_done_x112) begin
      res_0_sum <= res_0_sum + score_0_x112;
      res_1_sum <= res_1_sum + score_1_x112;
      res_2_sum <= res_2_sum + score_2_x112;
      res_3_sum <= res_3_sum + score_3_x112;
      res_4_sum <= res_4_sum + score_4_x112;
      res_5_sum <= res_5_sum + score_5_x112;
      res_6_sum <= res_6_sum + score_6_x112;
      res_7_sum <= res_7_sum + score_7_x112;
      res_8_sum <= res_8_sum + score_8_x112;
      res_9_sum <= res_9_sum + score_9_x112;
   end
   else if(res_done_x113) begin
      res_0_sum <= res_0_sum + score_0_x113;
      res_1_sum <= res_1_sum + score_1_x113;
      res_2_sum <= res_2_sum + score_2_x113;
      res_3_sum <= res_3_sum + score_3_x113;
      res_4_sum <= res_4_sum + score_4_x113;
      res_5_sum <= res_5_sum + score_5_x113;
      res_6_sum <= res_6_sum + score_6_x113;
      res_7_sum <= res_7_sum + score_7_x113;
      res_8_sum <= res_8_sum + score_8_x113;
      res_9_sum <= res_9_sum + score_9_x113;
   end
   else if(res_done_x114) begin
      res_0_sum <= res_0_sum + score_0_x114;
      res_1_sum <= res_1_sum + score_1_x114;
      res_2_sum <= res_2_sum + score_2_x114;
      res_3_sum <= res_3_sum + score_3_x114;
      res_4_sum <= res_4_sum + score_4_x114;
      res_5_sum <= res_5_sum + score_5_x114;
      res_6_sum <= res_6_sum + score_6_x114;
      res_7_sum <= res_7_sum + score_7_x114;
      res_8_sum <= res_8_sum + score_8_x114;
      res_9_sum <= res_9_sum + score_9_x114;
   end
   else if(res_done_x115) begin
      res_0_sum <= res_0_sum + score_0_x115;
      res_1_sum <= res_1_sum + score_1_x115;
      res_2_sum <= res_2_sum + score_2_x115;
      res_3_sum <= res_3_sum + score_3_x115;
      res_4_sum <= res_4_sum + score_4_x115;
      res_5_sum <= res_5_sum + score_5_x115;
      res_6_sum <= res_6_sum + score_6_x115;
      res_7_sum <= res_7_sum + score_7_x115;
      res_8_sum <= res_8_sum + score_8_x115;
      res_9_sum <= res_9_sum + score_9_x115;
   end
   else if(res_done_x116) begin
      res_0_sum <= res_0_sum + score_0_x116;
      res_1_sum <= res_1_sum + score_1_x116;
      res_2_sum <= res_2_sum + score_2_x116;
      res_3_sum <= res_3_sum + score_3_x116;
      res_4_sum <= res_4_sum + score_4_x116;
      res_5_sum <= res_5_sum + score_5_x116;
      res_6_sum <= res_6_sum + score_6_x116;
      res_7_sum <= res_7_sum + score_7_x116;
      res_8_sum <= res_8_sum + score_8_x116;
      res_9_sum <= res_9_sum + score_9_x116;
   end
   else if(res_done_x117) begin
      res_0_sum <= res_0_sum + score_0_x117;
      res_1_sum <= res_1_sum + score_1_x117;
      res_2_sum <= res_2_sum + score_2_x117;
      res_3_sum <= res_3_sum + score_3_x117;
      res_4_sum <= res_4_sum + score_4_x117;
      res_5_sum <= res_5_sum + score_5_x117;
      res_6_sum <= res_6_sum + score_6_x117;
      res_7_sum <= res_7_sum + score_7_x117;
      res_8_sum <= res_8_sum + score_8_x117;
      res_9_sum <= res_9_sum + score_9_x117;
   end
   else if(res_done_x118) begin
      res_0_sum <= res_0_sum + score_0_x118;
      res_1_sum <= res_1_sum + score_1_x118;
      res_2_sum <= res_2_sum + score_2_x118;
      res_3_sum <= res_3_sum + score_3_x118;
      res_4_sum <= res_4_sum + score_4_x118;
      res_5_sum <= res_5_sum + score_5_x118;
      res_6_sum <= res_6_sum + score_6_x118;
      res_7_sum <= res_7_sum + score_7_x118;
      res_8_sum <= res_8_sum + score_8_x118;
      res_9_sum <= res_9_sum + score_9_x118;
   end
   else if(res_done_x119) begin
      res_0_sum <= res_0_sum + score_0_x119;
      res_1_sum <= res_1_sum + score_1_x119;
      res_2_sum <= res_2_sum + score_2_x119;
      res_3_sum <= res_3_sum + score_3_x119;
      res_4_sum <= res_4_sum + score_4_x119;
      res_5_sum <= res_5_sum + score_5_x119;
      res_6_sum <= res_6_sum + score_6_x119;
      res_7_sum <= res_7_sum + score_7_x119;
      res_8_sum <= res_8_sum + score_8_x119;
      res_9_sum <= res_9_sum + score_9_x119;
   end
   else if(res_done_x120) begin
      res_0_sum <= res_0_sum + score_0_x120;
      res_1_sum <= res_1_sum + score_1_x120;
      res_2_sum <= res_2_sum + score_2_x120;
      res_3_sum <= res_3_sum + score_3_x120;
      res_4_sum <= res_4_sum + score_4_x120;
      res_5_sum <= res_5_sum + score_5_x120;
      res_6_sum <= res_6_sum + score_6_x120;
      res_7_sum <= res_7_sum + score_7_x120;
      res_8_sum <= res_8_sum + score_8_x120;
      res_9_sum <= res_9_sum + score_9_x120;
   end
   else if(res_done_x121) begin
      res_0_sum <= res_0_sum + score_0_x121;
      res_1_sum <= res_1_sum + score_1_x121;
      res_2_sum <= res_2_sum + score_2_x121;
      res_3_sum <= res_3_sum + score_3_x121;
      res_4_sum <= res_4_sum + score_4_x121;
      res_5_sum <= res_5_sum + score_5_x121;
      res_6_sum <= res_6_sum + score_6_x121;
      res_7_sum <= res_7_sum + score_7_x121;
      res_8_sum <= res_8_sum + score_8_x121;
      res_9_sum <= res_9_sum + score_9_x121;
   end
   else if(res_done_x122) begin
      res_0_sum <= res_0_sum + score_0_x122;
      res_1_sum <= res_1_sum + score_1_x122;
      res_2_sum <= res_2_sum + score_2_x122;
      res_3_sum <= res_3_sum + score_3_x122;
      res_4_sum <= res_4_sum + score_4_x122;
      res_5_sum <= res_5_sum + score_5_x122;
      res_6_sum <= res_6_sum + score_6_x122;
      res_7_sum <= res_7_sum + score_7_x122;
      res_8_sum <= res_8_sum + score_8_x122;
      res_9_sum <= res_9_sum + score_9_x122;
   end
   else if(res_done_x123) begin
      res_0_sum <= res_0_sum + score_0_x123;
      res_1_sum <= res_1_sum + score_1_x123;
      res_2_sum <= res_2_sum + score_2_x123;
      res_3_sum <= res_3_sum + score_3_x123;
      res_4_sum <= res_4_sum + score_4_x123;
      res_5_sum <= res_5_sum + score_5_x123;
      res_6_sum <= res_6_sum + score_6_x123;
      res_7_sum <= res_7_sum + score_7_x123;
      res_8_sum <= res_8_sum + score_8_x123;
      res_9_sum <= res_9_sum + score_9_x123;
   end
   else if(res_done_x124) begin
      res_0_sum <= res_0_sum + score_0_x124;
      res_1_sum <= res_1_sum + score_1_x124;
      res_2_sum <= res_2_sum + score_2_x124;
      res_3_sum <= res_3_sum + score_3_x124;
      res_4_sum <= res_4_sum + score_4_x124;
      res_5_sum <= res_5_sum + score_5_x124;
      res_6_sum <= res_6_sum + score_6_x124;
      res_7_sum <= res_7_sum + score_7_x124;
      res_8_sum <= res_8_sum + score_8_x124;
      res_9_sum <= res_9_sum + score_9_x124;
   end
   else if(res_done_x125) begin
      res_0_sum <= res_0_sum + score_0_x125;
      res_1_sum <= res_1_sum + score_1_x125;
      res_2_sum <= res_2_sum + score_2_x125;
      res_3_sum <= res_3_sum + score_3_x125;
      res_4_sum <= res_4_sum + score_4_x125;
      res_5_sum <= res_5_sum + score_5_x125;
      res_6_sum <= res_6_sum + score_6_x125;
      res_7_sum <= res_7_sum + score_7_x125;
      res_8_sum <= res_8_sum + score_8_x125;
      res_9_sum <= res_9_sum + score_9_x125;
   end
   else if(res_done_x126) begin
      res_0_sum <= res_0_sum + score_0_x126;
      res_1_sum <= res_1_sum + score_1_x126;
      res_2_sum <= res_2_sum + score_2_x126;
      res_3_sum <= res_3_sum + score_3_x126;
      res_4_sum <= res_4_sum + score_4_x126;
      res_5_sum <= res_5_sum + score_5_x126;
      res_6_sum <= res_6_sum + score_6_x126;
      res_7_sum <= res_7_sum + score_7_x126;
      res_8_sum <= res_8_sum + score_8_x126;
      res_9_sum <= res_9_sum + score_9_x126;
   end
   else if(res_done_x127) begin
      res_0_sum <= res_0_sum + score_0_x127;
      res_1_sum <= res_1_sum + score_1_x127;
      res_2_sum <= res_2_sum + score_2_x127;
      res_3_sum <= res_3_sum + score_3_x127;
      res_4_sum <= res_4_sum + score_4_x127;
      res_5_sum <= res_5_sum + score_5_x127;
      res_6_sum <= res_6_sum + score_6_x127;
      res_7_sum <= res_7_sum + score_7_x127;
      res_8_sum <= res_8_sum + score_8_x127;
      res_9_sum <= res_9_sum + score_9_x127;
   end
   else if(res_done_x128) begin
      res_0_sum <= res_0_sum + score_0_x128;
      res_1_sum <= res_1_sum + score_1_x128;
      res_2_sum <= res_2_sum + score_2_x128;
      res_3_sum <= res_3_sum + score_3_x128;
      res_4_sum <= res_4_sum + score_4_x128;
      res_5_sum <= res_5_sum + score_5_x128;
      res_6_sum <= res_6_sum + score_6_x128;
      res_7_sum <= res_7_sum + score_7_x128;
      res_8_sum <= res_8_sum + score_8_x128;
      res_9_sum <= res_9_sum + score_9_x128;
   end
   else if(res_done_x129) begin
      res_0_sum <= res_0_sum + score_0_x129;
      res_1_sum <= res_1_sum + score_1_x129;
      res_2_sum <= res_2_sum + score_2_x129;
      res_3_sum <= res_3_sum + score_3_x129;
      res_4_sum <= res_4_sum + score_4_x129;
      res_5_sum <= res_5_sum + score_5_x129;
      res_6_sum <= res_6_sum + score_6_x129;
      res_7_sum <= res_7_sum + score_7_x129;
      res_8_sum <= res_8_sum + score_8_x129;
      res_9_sum <= res_9_sum + score_9_x129;
   end
   else if(res_done_x130) begin
      res_0_sum <= res_0_sum + score_0_x130;
      res_1_sum <= res_1_sum + score_1_x130;
      res_2_sum <= res_2_sum + score_2_x130;
      res_3_sum <= res_3_sum + score_3_x130;
      res_4_sum <= res_4_sum + score_4_x130;
      res_5_sum <= res_5_sum + score_5_x130;
      res_6_sum <= res_6_sum + score_6_x130;
      res_7_sum <= res_7_sum + score_7_x130;
      res_8_sum <= res_8_sum + score_8_x130;
      res_9_sum <= res_9_sum + score_9_x130;
   end
   else if(res_done_x131) begin
      res_0_sum <= res_0_sum + score_0_x131;
      res_1_sum <= res_1_sum + score_1_x131;
      res_2_sum <= res_2_sum + score_2_x131;
      res_3_sum <= res_3_sum + score_3_x131;
      res_4_sum <= res_4_sum + score_4_x131;
      res_5_sum <= res_5_sum + score_5_x131;
      res_6_sum <= res_6_sum + score_6_x131;
      res_7_sum <= res_7_sum + score_7_x131;
      res_8_sum <= res_8_sum + score_8_x131;
      res_9_sum <= res_9_sum + score_9_x131;
   end
   else if(res_done_x132) begin
      res_0_sum <= res_0_sum + score_0_x132;
      res_1_sum <= res_1_sum + score_1_x132;
      res_2_sum <= res_2_sum + score_2_x132;
      res_3_sum <= res_3_sum + score_3_x132;
      res_4_sum <= res_4_sum + score_4_x132;
      res_5_sum <= res_5_sum + score_5_x132;
      res_6_sum <= res_6_sum + score_6_x132;
      res_7_sum <= res_7_sum + score_7_x132;
      res_8_sum <= res_8_sum + score_8_x132;
      res_9_sum <= res_9_sum + score_9_x132;
   end
   else if(res_done_x133) begin
      res_0_sum <= res_0_sum + score_0_x133;
      res_1_sum <= res_1_sum + score_1_x133;
      res_2_sum <= res_2_sum + score_2_x133;
      res_3_sum <= res_3_sum + score_3_x133;
      res_4_sum <= res_4_sum + score_4_x133;
      res_5_sum <= res_5_sum + score_5_x133;
      res_6_sum <= res_6_sum + score_6_x133;
      res_7_sum <= res_7_sum + score_7_x133;
      res_8_sum <= res_8_sum + score_8_x133;
      res_9_sum <= res_9_sum + score_9_x133;
   end
   else if(res_done_x134) begin
      res_0_sum <= res_0_sum + score_0_x134;
      res_1_sum <= res_1_sum + score_1_x134;
      res_2_sum <= res_2_sum + score_2_x134;
      res_3_sum <= res_3_sum + score_3_x134;
      res_4_sum <= res_4_sum + score_4_x134;
      res_5_sum <= res_5_sum + score_5_x134;
      res_6_sum <= res_6_sum + score_6_x134;
      res_7_sum <= res_7_sum + score_7_x134;
      res_8_sum <= res_8_sum + score_8_x134;
      res_9_sum <= res_9_sum + score_9_x134;
   end
   else if(res_done_x135) begin
      res_0_sum <= res_0_sum + score_0_x135;
      res_1_sum <= res_1_sum + score_1_x135;
      res_2_sum <= res_2_sum + score_2_x135;
      res_3_sum <= res_3_sum + score_3_x135;
      res_4_sum <= res_4_sum + score_4_x135;
      res_5_sum <= res_5_sum + score_5_x135;
      res_6_sum <= res_6_sum + score_6_x135;
      res_7_sum <= res_7_sum + score_7_x135;
      res_8_sum <= res_8_sum + score_8_x135;
      res_9_sum <= res_9_sum + score_9_x135;
   end
   else if(res_done_x136) begin
      res_0_sum <= res_0_sum + score_0_x136;
      res_1_sum <= res_1_sum + score_1_x136;
      res_2_sum <= res_2_sum + score_2_x136;
      res_3_sum <= res_3_sum + score_3_x136;
      res_4_sum <= res_4_sum + score_4_x136;
      res_5_sum <= res_5_sum + score_5_x136;
      res_6_sum <= res_6_sum + score_6_x136;
      res_7_sum <= res_7_sum + score_7_x136;
      res_8_sum <= res_8_sum + score_8_x136;
      res_9_sum <= res_9_sum + score_9_x136;
   end
   else if(res_done_x137) begin
      res_0_sum <= res_0_sum + score_0_x137;
      res_1_sum <= res_1_sum + score_1_x137;
      res_2_sum <= res_2_sum + score_2_x137;
      res_3_sum <= res_3_sum + score_3_x137;
      res_4_sum <= res_4_sum + score_4_x137;
      res_5_sum <= res_5_sum + score_5_x137;
      res_6_sum <= res_6_sum + score_6_x137;
      res_7_sum <= res_7_sum + score_7_x137;
      res_8_sum <= res_8_sum + score_8_x137;
      res_9_sum <= res_9_sum + score_9_x137;
   end
   else if(res_done_x138) begin
      res_0_sum <= res_0_sum + score_0_x138;
      res_1_sum <= res_1_sum + score_1_x138;
      res_2_sum <= res_2_sum + score_2_x138;
      res_3_sum <= res_3_sum + score_3_x138;
      res_4_sum <= res_4_sum + score_4_x138;
      res_5_sum <= res_5_sum + score_5_x138;
      res_6_sum <= res_6_sum + score_6_x138;
      res_7_sum <= res_7_sum + score_7_x138;
      res_8_sum <= res_8_sum + score_8_x138;
      res_9_sum <= res_9_sum + score_9_x138;
   end
   else if(res_done_x139) begin
      res_0_sum <= res_0_sum + score_0_x139;
      res_1_sum <= res_1_sum + score_1_x139;
      res_2_sum <= res_2_sum + score_2_x139;
      res_3_sum <= res_3_sum + score_3_x139;
      res_4_sum <= res_4_sum + score_4_x139;
      res_5_sum <= res_5_sum + score_5_x139;
      res_6_sum <= res_6_sum + score_6_x139;
      res_7_sum <= res_7_sum + score_7_x139;
      res_8_sum <= res_8_sum + score_8_x139;
      res_9_sum <= res_9_sum + score_9_x139;
   end
   else if(res_done_x140) begin
      res_0_sum <= res_0_sum + score_0_x140;
      res_1_sum <= res_1_sum + score_1_x140;
      res_2_sum <= res_2_sum + score_2_x140;
      res_3_sum <= res_3_sum + score_3_x140;
      res_4_sum <= res_4_sum + score_4_x140;
      res_5_sum <= res_5_sum + score_5_x140;
      res_6_sum <= res_6_sum + score_6_x140;
      res_7_sum <= res_7_sum + score_7_x140;
      res_8_sum <= res_8_sum + score_8_x140;
      res_9_sum <= res_9_sum + score_9_x140;
   end
   else if(res_done_x141) begin
      res_0_sum <= res_0_sum + score_0_x141;
      res_1_sum <= res_1_sum + score_1_x141;
      res_2_sum <= res_2_sum + score_2_x141;
      res_3_sum <= res_3_sum + score_3_x141;
      res_4_sum <= res_4_sum + score_4_x141;
      res_5_sum <= res_5_sum + score_5_x141;
      res_6_sum <= res_6_sum + score_6_x141;
      res_7_sum <= res_7_sum + score_7_x141;
      res_8_sum <= res_8_sum + score_8_x141;
      res_9_sum <= res_9_sum + score_9_x141;
   end
   else if(res_done_x142) begin
      res_0_sum <= res_0_sum + score_0_x142;
      res_1_sum <= res_1_sum + score_1_x142;
      res_2_sum <= res_2_sum + score_2_x142;
      res_3_sum <= res_3_sum + score_3_x142;
      res_4_sum <= res_4_sum + score_4_x142;
      res_5_sum <= res_5_sum + score_5_x142;
      res_6_sum <= res_6_sum + score_6_x142;
      res_7_sum <= res_7_sum + score_7_x142;
      res_8_sum <= res_8_sum + score_8_x142;
      res_9_sum <= res_9_sum + score_9_x142;
   end
   else if(res_done_x143) begin
      res_0_sum <= res_0_sum + score_0_x143;
      res_1_sum <= res_1_sum + score_1_x143;
      res_2_sum <= res_2_sum + score_2_x143;
      res_3_sum <= res_3_sum + score_3_x143;
      res_4_sum <= res_4_sum + score_4_x143;
      res_5_sum <= res_5_sum + score_5_x143;
      res_6_sum <= res_6_sum + score_6_x143;
      res_7_sum <= res_7_sum + score_7_x143;
      res_8_sum <= res_8_sum + score_8_x143;
      res_9_sum <= res_9_sum + score_9_x143;
   end
   else if(res_done_x144) begin
      res_0_sum <= res_0_sum + score_0_x144;
      res_1_sum <= res_1_sum + score_1_x144;
      res_2_sum <= res_2_sum + score_2_x144;
      res_3_sum <= res_3_sum + score_3_x144;
      res_4_sum <= res_4_sum + score_4_x144;
      res_5_sum <= res_5_sum + score_5_x144;
      res_6_sum <= res_6_sum + score_6_x144;
      res_7_sum <= res_7_sum + score_7_x144;
      res_8_sum <= res_8_sum + score_8_x144;
      res_9_sum <= res_9_sum + score_9_x144;
   end
   else if(res_done_x145) begin
      res_0_sum <= res_0_sum + score_0_x145;
      res_1_sum <= res_1_sum + score_1_x145;
      res_2_sum <= res_2_sum + score_2_x145;
      res_3_sum <= res_3_sum + score_3_x145;
      res_4_sum <= res_4_sum + score_4_x145;
      res_5_sum <= res_5_sum + score_5_x145;
      res_6_sum <= res_6_sum + score_6_x145;
      res_7_sum <= res_7_sum + score_7_x145;
      res_8_sum <= res_8_sum + score_8_x145;
      res_9_sum <= res_9_sum + score_9_x145;
   end
   else if(res_done_x146) begin
      res_0_sum <= res_0_sum + score_0_x146;
      res_1_sum <= res_1_sum + score_1_x146;
      res_2_sum <= res_2_sum + score_2_x146;
      res_3_sum <= res_3_sum + score_3_x146;
      res_4_sum <= res_4_sum + score_4_x146;
      res_5_sum <= res_5_sum + score_5_x146;
      res_6_sum <= res_6_sum + score_6_x146;
      res_7_sum <= res_7_sum + score_7_x146;
      res_8_sum <= res_8_sum + score_8_x146;
      res_9_sum <= res_9_sum + score_9_x146;
   end
   else if(res_done_x147) begin
      res_0_sum <= res_0_sum + score_0_x147;
      res_1_sum <= res_1_sum + score_1_x147;
      res_2_sum <= res_2_sum + score_2_x147;
      res_3_sum <= res_3_sum + score_3_x147;
      res_4_sum <= res_4_sum + score_4_x147;
      res_5_sum <= res_5_sum + score_5_x147;
      res_6_sum <= res_6_sum + score_6_x147;
      res_7_sum <= res_7_sum + score_7_x147;
      res_8_sum <= res_8_sum + score_8_x147;
      res_9_sum <= res_9_sum + score_9_x147;
   end
   else if(res_done_x148) begin
      res_0_sum <= res_0_sum + score_0_x148;
      res_1_sum <= res_1_sum + score_1_x148;
      res_2_sum <= res_2_sum + score_2_x148;
      res_3_sum <= res_3_sum + score_3_x148;
      res_4_sum <= res_4_sum + score_4_x148;
      res_5_sum <= res_5_sum + score_5_x148;
      res_6_sum <= res_6_sum + score_6_x148;
      res_7_sum <= res_7_sum + score_7_x148;
      res_8_sum <= res_8_sum + score_8_x148;
      res_9_sum <= res_9_sum + score_9_x148;
   end
   else if(res_done_x149) begin
      res_0_sum <= res_0_sum + score_0_x149;
      res_1_sum <= res_1_sum + score_1_x149;
      res_2_sum <= res_2_sum + score_2_x149;
      res_3_sum <= res_3_sum + score_3_x149;
      res_4_sum <= res_4_sum + score_4_x149;
      res_5_sum <= res_5_sum + score_5_x149;
      res_6_sum <= res_6_sum + score_6_x149;
      res_7_sum <= res_7_sum + score_7_x149;
      res_8_sum <= res_8_sum + score_8_x149;
      res_9_sum <= res_9_sum + score_9_x149;
   end
   else if(res_done_x150) begin
      res_0_sum <= res_0_sum + score_0_x150;
      res_1_sum <= res_1_sum + score_1_x150;
      res_2_sum <= res_2_sum + score_2_x150;
      res_3_sum <= res_3_sum + score_3_x150;
      res_4_sum <= res_4_sum + score_4_x150;
      res_5_sum <= res_5_sum + score_5_x150;
      res_6_sum <= res_6_sum + score_6_x150;
      res_7_sum <= res_7_sum + score_7_x150;
      res_8_sum <= res_8_sum + score_8_x150;
      res_9_sum <= res_9_sum + score_9_x150;
   end
   else if(res_done_x151) begin
      res_0_sum <= res_0_sum + score_0_x151;
      res_1_sum <= res_1_sum + score_1_x151;
      res_2_sum <= res_2_sum + score_2_x151;
      res_3_sum <= res_3_sum + score_3_x151;
      res_4_sum <= res_4_sum + score_4_x151;
      res_5_sum <= res_5_sum + score_5_x151;
      res_6_sum <= res_6_sum + score_6_x151;
      res_7_sum <= res_7_sum + score_7_x151;
      res_8_sum <= res_8_sum + score_8_x151;
      res_9_sum <= res_9_sum + score_9_x151;
   end
   else if(res_done_x152) begin
      res_0_sum <= res_0_sum + score_0_x152;
      res_1_sum <= res_1_sum + score_1_x152;
      res_2_sum <= res_2_sum + score_2_x152;
      res_3_sum <= res_3_sum + score_3_x152;
      res_4_sum <= res_4_sum + score_4_x152;
      res_5_sum <= res_5_sum + score_5_x152;
      res_6_sum <= res_6_sum + score_6_x152;
      res_7_sum <= res_7_sum + score_7_x152;
      res_8_sum <= res_8_sum + score_8_x152;
      res_9_sum <= res_9_sum + score_9_x152;
   end
   else if(res_done_x153) begin
      res_0_sum <= res_0_sum + score_0_x153;
      res_1_sum <= res_1_sum + score_1_x153;
      res_2_sum <= res_2_sum + score_2_x153;
      res_3_sum <= res_3_sum + score_3_x153;
      res_4_sum <= res_4_sum + score_4_x153;
      res_5_sum <= res_5_sum + score_5_x153;
      res_6_sum <= res_6_sum + score_6_x153;
      res_7_sum <= res_7_sum + score_7_x153;
      res_8_sum <= res_8_sum + score_8_x153;
      res_9_sum <= res_9_sum + score_9_x153;
   end
   else if(res_done_x154) begin
      res_0_sum <= res_0_sum + score_0_x154;
      res_1_sum <= res_1_sum + score_1_x154;
      res_2_sum <= res_2_sum + score_2_x154;
      res_3_sum <= res_3_sum + score_3_x154;
      res_4_sum <= res_4_sum + score_4_x154;
      res_5_sum <= res_5_sum + score_5_x154;
      res_6_sum <= res_6_sum + score_6_x154;
      res_7_sum <= res_7_sum + score_7_x154;
      res_8_sum <= res_8_sum + score_8_x154;
      res_9_sum <= res_9_sum + score_9_x154;
   end
   else if(res_done_x155) begin
      res_0_sum <= res_0_sum + score_0_x155;
      res_1_sum <= res_1_sum + score_1_x155;
      res_2_sum <= res_2_sum + score_2_x155;
      res_3_sum <= res_3_sum + score_3_x155;
      res_4_sum <= res_4_sum + score_4_x155;
      res_5_sum <= res_5_sum + score_5_x155;
      res_6_sum <= res_6_sum + score_6_x155;
      res_7_sum <= res_7_sum + score_7_x155;
      res_8_sum <= res_8_sum + score_8_x155;
      res_9_sum <= res_9_sum + score_9_x155;
   end
   else if(res_done_x156) begin
      res_0_sum <= res_0_sum + score_0_x156;
      res_1_sum <= res_1_sum + score_1_x156;
      res_2_sum <= res_2_sum + score_2_x156;
      res_3_sum <= res_3_sum + score_3_x156;
      res_4_sum <= res_4_sum + score_4_x156;
      res_5_sum <= res_5_sum + score_5_x156;
      res_6_sum <= res_6_sum + score_6_x156;
      res_7_sum <= res_7_sum + score_7_x156;
      res_8_sum <= res_8_sum + score_8_x156;
      res_9_sum <= res_9_sum + score_9_x156;
   end
   else if(res_done_x157) begin
      res_0_sum <= res_0_sum + score_0_x157;
      res_1_sum <= res_1_sum + score_1_x157;
      res_2_sum <= res_2_sum + score_2_x157;
      res_3_sum <= res_3_sum + score_3_x157;
      res_4_sum <= res_4_sum + score_4_x157;
      res_5_sum <= res_5_sum + score_5_x157;
      res_6_sum <= res_6_sum + score_6_x157;
      res_7_sum <= res_7_sum + score_7_x157;
      res_8_sum <= res_8_sum + score_8_x157;
      res_9_sum <= res_9_sum + score_9_x157;
   end
   else if(res_done_x158) begin
      res_0_sum <= res_0_sum + score_0_x158;
      res_1_sum <= res_1_sum + score_1_x158;
      res_2_sum <= res_2_sum + score_2_x158;
      res_3_sum <= res_3_sum + score_3_x158;
      res_4_sum <= res_4_sum + score_4_x158;
      res_5_sum <= res_5_sum + score_5_x158;
      res_6_sum <= res_6_sum + score_6_x158;
      res_7_sum <= res_7_sum + score_7_x158;
      res_8_sum <= res_8_sum + score_8_x158;
      res_9_sum <= res_9_sum + score_9_x158;
   end
   else if(res_done_x159) begin
      res_0_sum <= res_0_sum + score_0_x159;
      res_1_sum <= res_1_sum + score_1_x159;
      res_2_sum <= res_2_sum + score_2_x159;
      res_3_sum <= res_3_sum + score_3_x159;
      res_4_sum <= res_4_sum + score_4_x159;
      res_5_sum <= res_5_sum + score_5_x159;
      res_6_sum <= res_6_sum + score_6_x159;
      res_7_sum <= res_7_sum + score_7_x159;
      res_8_sum <= res_8_sum + score_8_x159;
      res_9_sum <= res_9_sum + score_9_x159;
   end
   else if(res_done_x160) begin
      res_0_sum <= res_0_sum + score_0_x160;
      res_1_sum <= res_1_sum + score_1_x160;
      res_2_sum <= res_2_sum + score_2_x160;
      res_3_sum <= res_3_sum + score_3_x160;
      res_4_sum <= res_4_sum + score_4_x160;
      res_5_sum <= res_5_sum + score_5_x160;
      res_6_sum <= res_6_sum + score_6_x160;
      res_7_sum <= res_7_sum + score_7_x160;
      res_8_sum <= res_8_sum + score_8_x160;
      res_9_sum <= res_9_sum + score_9_x160;
   end
   else if(res_done_x161) begin
      res_0_sum <= res_0_sum + score_0_x161;
      res_1_sum <= res_1_sum + score_1_x161;
      res_2_sum <= res_2_sum + score_2_x161;
      res_3_sum <= res_3_sum + score_3_x161;
      res_4_sum <= res_4_sum + score_4_x161;
      res_5_sum <= res_5_sum + score_5_x161;
      res_6_sum <= res_6_sum + score_6_x161;
      res_7_sum <= res_7_sum + score_7_x161;
      res_8_sum <= res_8_sum + score_8_x161;
      res_9_sum <= res_9_sum + score_9_x161;
   end
   else if(res_done_x162) begin
      res_0_sum <= res_0_sum + score_0_x162;
      res_1_sum <= res_1_sum + score_1_x162;
      res_2_sum <= res_2_sum + score_2_x162;
      res_3_sum <= res_3_sum + score_3_x162;
      res_4_sum <= res_4_sum + score_4_x162;
      res_5_sum <= res_5_sum + score_5_x162;
      res_6_sum <= res_6_sum + score_6_x162;
      res_7_sum <= res_7_sum + score_7_x162;
      res_8_sum <= res_8_sum + score_8_x162;
      res_9_sum <= res_9_sum + score_9_x162;
   end
   else if(res_done_x163) begin
      res_0_sum <= res_0_sum + score_0_x163;
      res_1_sum <= res_1_sum + score_1_x163;
      res_2_sum <= res_2_sum + score_2_x163;
      res_3_sum <= res_3_sum + score_3_x163;
      res_4_sum <= res_4_sum + score_4_x163;
      res_5_sum <= res_5_sum + score_5_x163;
      res_6_sum <= res_6_sum + score_6_x163;
      res_7_sum <= res_7_sum + score_7_x163;
      res_8_sum <= res_8_sum + score_8_x163;
      res_9_sum <= res_9_sum + score_9_x163;
   end
   else if(res_done_x164) begin
      res_0_sum <= res_0_sum + score_0_x164;
      res_1_sum <= res_1_sum + score_1_x164;
      res_2_sum <= res_2_sum + score_2_x164;
      res_3_sum <= res_3_sum + score_3_x164;
      res_4_sum <= res_4_sum + score_4_x164;
      res_5_sum <= res_5_sum + score_5_x164;
      res_6_sum <= res_6_sum + score_6_x164;
      res_7_sum <= res_7_sum + score_7_x164;
      res_8_sum <= res_8_sum + score_8_x164;
      res_9_sum <= res_9_sum + score_9_x164;
   end
   else if(res_done_x165) begin
      res_0_sum <= res_0_sum + score_0_x165;
      res_1_sum <= res_1_sum + score_1_x165;
      res_2_sum <= res_2_sum + score_2_x165;
      res_3_sum <= res_3_sum + score_3_x165;
      res_4_sum <= res_4_sum + score_4_x165;
      res_5_sum <= res_5_sum + score_5_x165;
      res_6_sum <= res_6_sum + score_6_x165;
      res_7_sum <= res_7_sum + score_7_x165;
      res_8_sum <= res_8_sum + score_8_x165;
      res_9_sum <= res_9_sum + score_9_x165;
   end
   else if(res_done_x166) begin
      res_0_sum <= res_0_sum + score_0_x166;
      res_1_sum <= res_1_sum + score_1_x166;
      res_2_sum <= res_2_sum + score_2_x166;
      res_3_sum <= res_3_sum + score_3_x166;
      res_4_sum <= res_4_sum + score_4_x166;
      res_5_sum <= res_5_sum + score_5_x166;
      res_6_sum <= res_6_sum + score_6_x166;
      res_7_sum <= res_7_sum + score_7_x166;
      res_8_sum <= res_8_sum + score_8_x166;
      res_9_sum <= res_9_sum + score_9_x166;
   end
   else if(res_done_x167) begin
      res_0_sum <= res_0_sum + score_0_x167;
      res_1_sum <= res_1_sum + score_1_x167;
      res_2_sum <= res_2_sum + score_2_x167;
      res_3_sum <= res_3_sum + score_3_x167;
      res_4_sum <= res_4_sum + score_4_x167;
      res_5_sum <= res_5_sum + score_5_x167;
      res_6_sum <= res_6_sum + score_6_x167;
      res_7_sum <= res_7_sum + score_7_x167;
      res_8_sum <= res_8_sum + score_8_x167;
      res_9_sum <= res_9_sum + score_9_x167;
   end
   else if(res_done_x168) begin
      res_0_sum <= res_0_sum + score_0_x168;
      res_1_sum <= res_1_sum + score_1_x168;
      res_2_sum <= res_2_sum + score_2_x168;
      res_3_sum <= res_3_sum + score_3_x168;
      res_4_sum <= res_4_sum + score_4_x168;
      res_5_sum <= res_5_sum + score_5_x168;
      res_6_sum <= res_6_sum + score_6_x168;
      res_7_sum <= res_7_sum + score_7_x168;
      res_8_sum <= res_8_sum + score_8_x168;
      res_9_sum <= res_9_sum + score_9_x168;
   end
   else if(res_done_x169) begin
      res_0_sum <= res_0_sum + score_0_x169;
      res_1_sum <= res_1_sum + score_1_x169;
      res_2_sum <= res_2_sum + score_2_x169;
      res_3_sum <= res_3_sum + score_3_x169;
      res_4_sum <= res_4_sum + score_4_x169;
      res_5_sum <= res_5_sum + score_5_x169;
      res_6_sum <= res_6_sum + score_6_x169;
      res_7_sum <= res_7_sum + score_7_x169;
      res_8_sum <= res_8_sum + score_8_x169;
      res_9_sum <= res_9_sum + score_9_x169;
   end
   else if(res_done_x170) begin
      res_0_sum <= res_0_sum + score_0_x170;
      res_1_sum <= res_1_sum + score_1_x170;
      res_2_sum <= res_2_sum + score_2_x170;
      res_3_sum <= res_3_sum + score_3_x170;
      res_4_sum <= res_4_sum + score_4_x170;
      res_5_sum <= res_5_sum + score_5_x170;
      res_6_sum <= res_6_sum + score_6_x170;
      res_7_sum <= res_7_sum + score_7_x170;
      res_8_sum <= res_8_sum + score_8_x170;
      res_9_sum <= res_9_sum + score_9_x170;
   end
   else if(res_done_x171) begin
      res_0_sum <= res_0_sum + score_0_x171;
      res_1_sum <= res_1_sum + score_1_x171;
      res_2_sum <= res_2_sum + score_2_x171;
      res_3_sum <= res_3_sum + score_3_x171;
      res_4_sum <= res_4_sum + score_4_x171;
      res_5_sum <= res_5_sum + score_5_x171;
      res_6_sum <= res_6_sum + score_6_x171;
      res_7_sum <= res_7_sum + score_7_x171;
      res_8_sum <= res_8_sum + score_8_x171;
      res_9_sum <= res_9_sum + score_9_x171;
   end
   else if(res_done_x172) begin
      res_0_sum <= res_0_sum + score_0_x172;
      res_1_sum <= res_1_sum + score_1_x172;
      res_2_sum <= res_2_sum + score_2_x172;
      res_3_sum <= res_3_sum + score_3_x172;
      res_4_sum <= res_4_sum + score_4_x172;
      res_5_sum <= res_5_sum + score_5_x172;
      res_6_sum <= res_6_sum + score_6_x172;
      res_7_sum <= res_7_sum + score_7_x172;
      res_8_sum <= res_8_sum + score_8_x172;
      res_9_sum <= res_9_sum + score_9_x172;
   end
   else if(res_done_x173) begin
      res_0_sum <= res_0_sum + score_0_x173;
      res_1_sum <= res_1_sum + score_1_x173;
      res_2_sum <= res_2_sum + score_2_x173;
      res_3_sum <= res_3_sum + score_3_x173;
      res_4_sum <= res_4_sum + score_4_x173;
      res_5_sum <= res_5_sum + score_5_x173;
      res_6_sum <= res_6_sum + score_6_x173;
      res_7_sum <= res_7_sum + score_7_x173;
      res_8_sum <= res_8_sum + score_8_x173;
      res_9_sum <= res_9_sum + score_9_x173;
   end
   else if(res_done_x174) begin
      res_0_sum <= res_0_sum + score_0_x174;
      res_1_sum <= res_1_sum + score_1_x174;
      res_2_sum <= res_2_sum + score_2_x174;
      res_3_sum <= res_3_sum + score_3_x174;
      res_4_sum <= res_4_sum + score_4_x174;
      res_5_sum <= res_5_sum + score_5_x174;
      res_6_sum <= res_6_sum + score_6_x174;
      res_7_sum <= res_7_sum + score_7_x174;
      res_8_sum <= res_8_sum + score_8_x174;
      res_9_sum <= res_9_sum + score_9_x174;
   end
   else if(res_done_x175) begin
      res_0_sum <= res_0_sum + score_0_x175;
      res_1_sum <= res_1_sum + score_1_x175;
      res_2_sum <= res_2_sum + score_2_x175;
      res_3_sum <= res_3_sum + score_3_x175;
      res_4_sum <= res_4_sum + score_4_x175;
      res_5_sum <= res_5_sum + score_5_x175;
      res_6_sum <= res_6_sum + score_6_x175;
      res_7_sum <= res_7_sum + score_7_x175;
      res_8_sum <= res_8_sum + score_8_x175;
      res_9_sum <= res_9_sum + score_9_x175;
   end
   else if(res_done_x176) begin
      res_0_sum <= res_0_sum + score_0_x176;
      res_1_sum <= res_1_sum + score_1_x176;
      res_2_sum <= res_2_sum + score_2_x176;
      res_3_sum <= res_3_sum + score_3_x176;
      res_4_sum <= res_4_sum + score_4_x176;
      res_5_sum <= res_5_sum + score_5_x176;
      res_6_sum <= res_6_sum + score_6_x176;
      res_7_sum <= res_7_sum + score_7_x176;
      res_8_sum <= res_8_sum + score_8_x176;
      res_9_sum <= res_9_sum + score_9_x176;
   end
   else if(res_done_x177) begin
      res_0_sum <= res_0_sum + score_0_x177;
      res_1_sum <= res_1_sum + score_1_x177;
      res_2_sum <= res_2_sum + score_2_x177;
      res_3_sum <= res_3_sum + score_3_x177;
      res_4_sum <= res_4_sum + score_4_x177;
      res_5_sum <= res_5_sum + score_5_x177;
      res_6_sum <= res_6_sum + score_6_x177;
      res_7_sum <= res_7_sum + score_7_x177;
      res_8_sum <= res_8_sum + score_8_x177;
      res_9_sum <= res_9_sum + score_9_x177;
   end
   else if(res_done_x178) begin
      res_0_sum <= res_0_sum + score_0_x178;
      res_1_sum <= res_1_sum + score_1_x178;
      res_2_sum <= res_2_sum + score_2_x178;
      res_3_sum <= res_3_sum + score_3_x178;
      res_4_sum <= res_4_sum + score_4_x178;
      res_5_sum <= res_5_sum + score_5_x178;
      res_6_sum <= res_6_sum + score_6_x178;
      res_7_sum <= res_7_sum + score_7_x178;
      res_8_sum <= res_8_sum + score_8_x178;
      res_9_sum <= res_9_sum + score_9_x178;
   end
   else if(res_done_x179) begin
      res_0_sum <= res_0_sum + score_0_x179;
      res_1_sum <= res_1_sum + score_1_x179;
      res_2_sum <= res_2_sum + score_2_x179;
      res_3_sum <= res_3_sum + score_3_x179;
      res_4_sum <= res_4_sum + score_4_x179;
      res_5_sum <= res_5_sum + score_5_x179;
      res_6_sum <= res_6_sum + score_6_x179;
      res_7_sum <= res_7_sum + score_7_x179;
      res_8_sum <= res_8_sum + score_8_x179;
      res_9_sum <= res_9_sum + score_9_x179;
   end
   else if(res_done_x180) begin
      res_0_sum <= res_0_sum + score_0_x180;
      res_1_sum <= res_1_sum + score_1_x180;
      res_2_sum <= res_2_sum + score_2_x180;
      res_3_sum <= res_3_sum + score_3_x180;
      res_4_sum <= res_4_sum + score_4_x180;
      res_5_sum <= res_5_sum + score_5_x180;
      res_6_sum <= res_6_sum + score_6_x180;
      res_7_sum <= res_7_sum + score_7_x180;
      res_8_sum <= res_8_sum + score_8_x180;
      res_9_sum <= res_9_sum + score_9_x180;
   end
   else if(res_done_x181) begin
      res_0_sum <= res_0_sum + score_0_x181;
      res_1_sum <= res_1_sum + score_1_x181;
      res_2_sum <= res_2_sum + score_2_x181;
      res_3_sum <= res_3_sum + score_3_x181;
      res_4_sum <= res_4_sum + score_4_x181;
      res_5_sum <= res_5_sum + score_5_x181;
      res_6_sum <= res_6_sum + score_6_x181;
      res_7_sum <= res_7_sum + score_7_x181;
      res_8_sum <= res_8_sum + score_8_x181;
      res_9_sum <= res_9_sum + score_9_x181;
   end
   else if(res_done_x182) begin
      res_0_sum <= res_0_sum + score_0_x182;
      res_1_sum <= res_1_sum + score_1_x182;
      res_2_sum <= res_2_sum + score_2_x182;
      res_3_sum <= res_3_sum + score_3_x182;
      res_4_sum <= res_4_sum + score_4_x182;
      res_5_sum <= res_5_sum + score_5_x182;
      res_6_sum <= res_6_sum + score_6_x182;
      res_7_sum <= res_7_sum + score_7_x182;
      res_8_sum <= res_8_sum + score_8_x182;
      res_9_sum <= res_9_sum + score_9_x182;
   end
   else if(res_done_x183) begin
      res_0_sum <= res_0_sum + score_0_x183;
      res_1_sum <= res_1_sum + score_1_x183;
      res_2_sum <= res_2_sum + score_2_x183;
      res_3_sum <= res_3_sum + score_3_x183;
      res_4_sum <= res_4_sum + score_4_x183;
      res_5_sum <= res_5_sum + score_5_x183;
      res_6_sum <= res_6_sum + score_6_x183;
      res_7_sum <= res_7_sum + score_7_x183;
      res_8_sum <= res_8_sum + score_8_x183;
      res_9_sum <= res_9_sum + score_9_x183;
   end
   else if(res_done_x184) begin
      res_0_sum <= res_0_sum + score_0_x184;
      res_1_sum <= res_1_sum + score_1_x184;
      res_2_sum <= res_2_sum + score_2_x184;
      res_3_sum <= res_3_sum + score_3_x184;
      res_4_sum <= res_4_sum + score_4_x184;
      res_5_sum <= res_5_sum + score_5_x184;
      res_6_sum <= res_6_sum + score_6_x184;
      res_7_sum <= res_7_sum + score_7_x184;
      res_8_sum <= res_8_sum + score_8_x184;
      res_9_sum <= res_9_sum + score_9_x184;
   end
   else if(res_done_x185) begin
      res_0_sum <= res_0_sum + score_0_x185;
      res_1_sum <= res_1_sum + score_1_x185;
      res_2_sum <= res_2_sum + score_2_x185;
      res_3_sum <= res_3_sum + score_3_x185;
      res_4_sum <= res_4_sum + score_4_x185;
      res_5_sum <= res_5_sum + score_5_x185;
      res_6_sum <= res_6_sum + score_6_x185;
      res_7_sum <= res_7_sum + score_7_x185;
      res_8_sum <= res_8_sum + score_8_x185;
      res_9_sum <= res_9_sum + score_9_x185;
   end
   else if(res_done_x186) begin
      res_0_sum <= res_0_sum + score_0_x186;
      res_1_sum <= res_1_sum + score_1_x186;
      res_2_sum <= res_2_sum + score_2_x186;
      res_3_sum <= res_3_sum + score_3_x186;
      res_4_sum <= res_4_sum + score_4_x186;
      res_5_sum <= res_5_sum + score_5_x186;
      res_6_sum <= res_6_sum + score_6_x186;
      res_7_sum <= res_7_sum + score_7_x186;
      res_8_sum <= res_8_sum + score_8_x186;
      res_9_sum <= res_9_sum + score_9_x186;
   end
   else if(res_done_x187) begin
      res_0_sum <= res_0_sum + score_0_x187;
      res_1_sum <= res_1_sum + score_1_x187;
      res_2_sum <= res_2_sum + score_2_x187;
      res_3_sum <= res_3_sum + score_3_x187;
      res_4_sum <= res_4_sum + score_4_x187;
      res_5_sum <= res_5_sum + score_5_x187;
      res_6_sum <= res_6_sum + score_6_x187;
      res_7_sum <= res_7_sum + score_7_x187;
      res_8_sum <= res_8_sum + score_8_x187;
      res_9_sum <= res_9_sum + score_9_x187;
   end
   else if(res_done_x188) begin
      res_0_sum <= res_0_sum + score_0_x188;
      res_1_sum <= res_1_sum + score_1_x188;
      res_2_sum <= res_2_sum + score_2_x188;
      res_3_sum <= res_3_sum + score_3_x188;
      res_4_sum <= res_4_sum + score_4_x188;
      res_5_sum <= res_5_sum + score_5_x188;
      res_6_sum <= res_6_sum + score_6_x188;
      res_7_sum <= res_7_sum + score_7_x188;
      res_8_sum <= res_8_sum + score_8_x188;
      res_9_sum <= res_9_sum + score_9_x188;
   end
   else if(res_done_x189) begin
      res_0_sum <= res_0_sum + score_0_x189;
      res_1_sum <= res_1_sum + score_1_x189;
      res_2_sum <= res_2_sum + score_2_x189;
      res_3_sum <= res_3_sum + score_3_x189;
      res_4_sum <= res_4_sum + score_4_x189;
      res_5_sum <= res_5_sum + score_5_x189;
      res_6_sum <= res_6_sum + score_6_x189;
      res_7_sum <= res_7_sum + score_7_x189;
      res_8_sum <= res_8_sum + score_8_x189;
      res_9_sum <= res_9_sum + score_9_x189;
   end
   else if(res_done_x190) begin
      res_0_sum <= res_0_sum + score_0_x190;
      res_1_sum <= res_1_sum + score_1_x190;
      res_2_sum <= res_2_sum + score_2_x190;
      res_3_sum <= res_3_sum + score_3_x190;
      res_4_sum <= res_4_sum + score_4_x190;
      res_5_sum <= res_5_sum + score_5_x190;
      res_6_sum <= res_6_sum + score_6_x190;
      res_7_sum <= res_7_sum + score_7_x190;
      res_8_sum <= res_8_sum + score_8_x190;
      res_9_sum <= res_9_sum + score_9_x190;
   end
   else if(res_done_x191) begin
      res_0_sum <= res_0_sum + score_0_x191;
      res_1_sum <= res_1_sum + score_1_x191;
      res_2_sum <= res_2_sum + score_2_x191;
      res_3_sum <= res_3_sum + score_3_x191;
      res_4_sum <= res_4_sum + score_4_x191;
      res_5_sum <= res_5_sum + score_5_x191;
      res_6_sum <= res_6_sum + score_6_x191;
      res_7_sum <= res_7_sum + score_7_x191;
      res_8_sum <= res_8_sum + score_8_x191;
      res_9_sum <= res_9_sum + score_9_x191;
   end
   else if(res_done_x192) begin
      res_0_sum <= res_0_sum + score_0_x192;
      res_1_sum <= res_1_sum + score_1_x192;
      res_2_sum <= res_2_sum + score_2_x192;
      res_3_sum <= res_3_sum + score_3_x192;
      res_4_sum <= res_4_sum + score_4_x192;
      res_5_sum <= res_5_sum + score_5_x192;
      res_6_sum <= res_6_sum + score_6_x192;
      res_7_sum <= res_7_sum + score_7_x192;
      res_8_sum <= res_8_sum + score_8_x192;
      res_9_sum <= res_9_sum + score_9_x192;
   end
   else if(res_done_x193) begin
      res_0_sum <= res_0_sum + score_0_x193;
      res_1_sum <= res_1_sum + score_1_x193;
      res_2_sum <= res_2_sum + score_2_x193;
      res_3_sum <= res_3_sum + score_3_x193;
      res_4_sum <= res_4_sum + score_4_x193;
      res_5_sum <= res_5_sum + score_5_x193;
      res_6_sum <= res_6_sum + score_6_x193;
      res_7_sum <= res_7_sum + score_7_x193;
      res_8_sum <= res_8_sum + score_8_x193;
      res_9_sum <= res_9_sum + score_9_x193;
   end
   else if(res_done_x194) begin
      res_0_sum <= res_0_sum + score_0_x194;
      res_1_sum <= res_1_sum + score_1_x194;
      res_2_sum <= res_2_sum + score_2_x194;
      res_3_sum <= res_3_sum + score_3_x194;
      res_4_sum <= res_4_sum + score_4_x194;
      res_5_sum <= res_5_sum + score_5_x194;
      res_6_sum <= res_6_sum + score_6_x194;
      res_7_sum <= res_7_sum + score_7_x194;
      res_8_sum <= res_8_sum + score_8_x194;
      res_9_sum <= res_9_sum + score_9_x194;
   end
   else if(res_done_x195) begin
      res_0_sum <= res_0_sum + score_0_x195;
      res_1_sum <= res_1_sum + score_1_x195;
      res_2_sum <= res_2_sum + score_2_x195;
      res_3_sum <= res_3_sum + score_3_x195;
      res_4_sum <= res_4_sum + score_4_x195;
      res_5_sum <= res_5_sum + score_5_x195;
      res_6_sum <= res_6_sum + score_6_x195;
      res_7_sum <= res_7_sum + score_7_x195;
      res_8_sum <= res_8_sum + score_8_x195;
      res_9_sum <= res_9_sum + score_9_x195;
   end
   else if(res_done_x196) begin
      res_0_sum <= res_0_sum + score_0_x196;
      res_1_sum <= res_1_sum + score_1_x196;
      res_2_sum <= res_2_sum + score_2_x196;
      res_3_sum <= res_3_sum + score_3_x196;
      res_4_sum <= res_4_sum + score_4_x196;
      res_5_sum <= res_5_sum + score_5_x196;
      res_6_sum <= res_6_sum + score_6_x196;
      res_7_sum <= res_7_sum + score_7_x196;
      res_8_sum <= res_8_sum + score_8_x196;
      res_9_sum <= res_9_sum + score_9_x196;
   end
   else if(res_done_x197) begin
      res_0_sum <= res_0_sum + score_0_x197;
      res_1_sum <= res_1_sum + score_1_x197;
      res_2_sum <= res_2_sum + score_2_x197;
      res_3_sum <= res_3_sum + score_3_x197;
      res_4_sum <= res_4_sum + score_4_x197;
      res_5_sum <= res_5_sum + score_5_x197;
      res_6_sum <= res_6_sum + score_6_x197;
      res_7_sum <= res_7_sum + score_7_x197;
      res_8_sum <= res_8_sum + score_8_x197;
      res_9_sum <= res_9_sum + score_9_x197;
   end
   else if(res_done_x198) begin
      res_0_sum <= res_0_sum + score_0_x198;
      res_1_sum <= res_1_sum + score_1_x198;
      res_2_sum <= res_2_sum + score_2_x198;
      res_3_sum <= res_3_sum + score_3_x198;
      res_4_sum <= res_4_sum + score_4_x198;
      res_5_sum <= res_5_sum + score_5_x198;
      res_6_sum <= res_6_sum + score_6_x198;
      res_7_sum <= res_7_sum + score_7_x198;
      res_8_sum <= res_8_sum + score_8_x198;
      res_9_sum <= res_9_sum + score_9_x198;
   end
   else if(res_done_x199) begin
      res_0_sum <= res_0_sum + score_0_x199;
      res_1_sum <= res_1_sum + score_1_x199;
      res_2_sum <= res_2_sum + score_2_x199;
      res_3_sum <= res_3_sum + score_3_x199;
      res_4_sum <= res_4_sum + score_4_x199;
      res_5_sum <= res_5_sum + score_5_x199;
      res_6_sum <= res_6_sum + score_6_x199;
      res_7_sum <= res_7_sum + score_7_x199;
      res_8_sum <= res_8_sum + score_8_x199;
      res_9_sum <= res_9_sum + score_9_x199;
   end
   else if(res_done_x200) begin
      res_0_sum <= res_0_sum + score_0_x200;
      res_1_sum <= res_1_sum + score_1_x200;
      res_2_sum <= res_2_sum + score_2_x200;
      res_3_sum <= res_3_sum + score_3_x200;
      res_4_sum <= res_4_sum + score_4_x200;
      res_5_sum <= res_5_sum + score_5_x200;
      res_6_sum <= res_6_sum + score_6_x200;
      res_7_sum <= res_7_sum + score_7_x200;
      res_8_sum <= res_8_sum + score_8_x200;
      res_9_sum <= res_9_sum + score_9_x200;
   end
   else if(res_done_x201) begin
      res_0_sum <= res_0_sum + score_0_x201;
      res_1_sum <= res_1_sum + score_1_x201;
      res_2_sum <= res_2_sum + score_2_x201;
      res_3_sum <= res_3_sum + score_3_x201;
      res_4_sum <= res_4_sum + score_4_x201;
      res_5_sum <= res_5_sum + score_5_x201;
      res_6_sum <= res_6_sum + score_6_x201;
      res_7_sum <= res_7_sum + score_7_x201;
      res_8_sum <= res_8_sum + score_8_x201;
      res_9_sum <= res_9_sum + score_9_x201;
   end
   else if(res_done_x202) begin
      res_0_sum <= res_0_sum + score_0_x202;
      res_1_sum <= res_1_sum + score_1_x202;
      res_2_sum <= res_2_sum + score_2_x202;
      res_3_sum <= res_3_sum + score_3_x202;
      res_4_sum <= res_4_sum + score_4_x202;
      res_5_sum <= res_5_sum + score_5_x202;
      res_6_sum <= res_6_sum + score_6_x202;
      res_7_sum <= res_7_sum + score_7_x202;
      res_8_sum <= res_8_sum + score_8_x202;
      res_9_sum <= res_9_sum + score_9_x202;
   end
   else if(res_done_x203) begin
      res_0_sum <= res_0_sum + score_0_x203;
      res_1_sum <= res_1_sum + score_1_x203;
      res_2_sum <= res_2_sum + score_2_x203;
      res_3_sum <= res_3_sum + score_3_x203;
      res_4_sum <= res_4_sum + score_4_x203;
      res_5_sum <= res_5_sum + score_5_x203;
      res_6_sum <= res_6_sum + score_6_x203;
      res_7_sum <= res_7_sum + score_7_x203;
      res_8_sum <= res_8_sum + score_8_x203;
      res_9_sum <= res_9_sum + score_9_x203;
   end
   else if(res_done_x204) begin
      res_0_sum <= res_0_sum + score_0_x204;
      res_1_sum <= res_1_sum + score_1_x204;
      res_2_sum <= res_2_sum + score_2_x204;
      res_3_sum <= res_3_sum + score_3_x204;
      res_4_sum <= res_4_sum + score_4_x204;
      res_5_sum <= res_5_sum + score_5_x204;
      res_6_sum <= res_6_sum + score_6_x204;
      res_7_sum <= res_7_sum + score_7_x204;
      res_8_sum <= res_8_sum + score_8_x204;
      res_9_sum <= res_9_sum + score_9_x204;
   end
   else if(res_done_x205) begin
      res_0_sum <= res_0_sum + score_0_x205;
      res_1_sum <= res_1_sum + score_1_x205;
      res_2_sum <= res_2_sum + score_2_x205;
      res_3_sum <= res_3_sum + score_3_x205;
      res_4_sum <= res_4_sum + score_4_x205;
      res_5_sum <= res_5_sum + score_5_x205;
      res_6_sum <= res_6_sum + score_6_x205;
      res_7_sum <= res_7_sum + score_7_x205;
      res_8_sum <= res_8_sum + score_8_x205;
      res_9_sum <= res_9_sum + score_9_x205;
   end
   else if(res_done_x206) begin
      res_0_sum <= res_0_sum + score_0_x206;
      res_1_sum <= res_1_sum + score_1_x206;
      res_2_sum <= res_2_sum + score_2_x206;
      res_3_sum <= res_3_sum + score_3_x206;
      res_4_sum <= res_4_sum + score_4_x206;
      res_5_sum <= res_5_sum + score_5_x206;
      res_6_sum <= res_6_sum + score_6_x206;
      res_7_sum <= res_7_sum + score_7_x206;
      res_8_sum <= res_8_sum + score_8_x206;
      res_9_sum <= res_9_sum + score_9_x206;
   end
   else if(res_done_x207) begin
      res_0_sum <= res_0_sum + score_0_x207;
      res_1_sum <= res_1_sum + score_1_x207;
      res_2_sum <= res_2_sum + score_2_x207;
      res_3_sum <= res_3_sum + score_3_x207;
      res_4_sum <= res_4_sum + score_4_x207;
      res_5_sum <= res_5_sum + score_5_x207;
      res_6_sum <= res_6_sum + score_6_x207;
      res_7_sum <= res_7_sum + score_7_x207;
      res_8_sum <= res_8_sum + score_8_x207;
      res_9_sum <= res_9_sum + score_9_x207;
   end
   else if(res_done_x208) begin
      res_0_sum <= res_0_sum + score_0_x208;
      res_1_sum <= res_1_sum + score_1_x208;
      res_2_sum <= res_2_sum + score_2_x208;
      res_3_sum <= res_3_sum + score_3_x208;
      res_4_sum <= res_4_sum + score_4_x208;
      res_5_sum <= res_5_sum + score_5_x208;
      res_6_sum <= res_6_sum + score_6_x208;
      res_7_sum <= res_7_sum + score_7_x208;
      res_8_sum <= res_8_sum + score_8_x208;
      res_9_sum <= res_9_sum + score_9_x208;
   end
   else if(res_done_x209) begin
      res_0_sum <= res_0_sum + score_0_x209;
      res_1_sum <= res_1_sum + score_1_x209;
      res_2_sum <= res_2_sum + score_2_x209;
      res_3_sum <= res_3_sum + score_3_x209;
      res_4_sum <= res_4_sum + score_4_x209;
      res_5_sum <= res_5_sum + score_5_x209;
      res_6_sum <= res_6_sum + score_6_x209;
      res_7_sum <= res_7_sum + score_7_x209;
      res_8_sum <= res_8_sum + score_8_x209;
      res_9_sum <= res_9_sum + score_9_x209;
   end
   else if(res_done_x210) begin
      res_0_sum <= res_0_sum + score_0_x210;
      res_1_sum <= res_1_sum + score_1_x210;
      res_2_sum <= res_2_sum + score_2_x210;
      res_3_sum <= res_3_sum + score_3_x210;
      res_4_sum <= res_4_sum + score_4_x210;
      res_5_sum <= res_5_sum + score_5_x210;
      res_6_sum <= res_6_sum + score_6_x210;
      res_7_sum <= res_7_sum + score_7_x210;
      res_8_sum <= res_8_sum + score_8_x210;
      res_9_sum <= res_9_sum + score_9_x210;
   end
   else if(res_done_x211) begin
      res_0_sum <= res_0_sum + score_0_x211;
      res_1_sum <= res_1_sum + score_1_x211;
      res_2_sum <= res_2_sum + score_2_x211;
      res_3_sum <= res_3_sum + score_3_x211;
      res_4_sum <= res_4_sum + score_4_x211;
      res_5_sum <= res_5_sum + score_5_x211;
      res_6_sum <= res_6_sum + score_6_x211;
      res_7_sum <= res_7_sum + score_7_x211;
      res_8_sum <= res_8_sum + score_8_x211;
      res_9_sum <= res_9_sum + score_9_x211;
   end
   else if(res_done_x212) begin
      res_0_sum <= res_0_sum + score_0_x212;
      res_1_sum <= res_1_sum + score_1_x212;
      res_2_sum <= res_2_sum + score_2_x212;
      res_3_sum <= res_3_sum + score_3_x212;
      res_4_sum <= res_4_sum + score_4_x212;
      res_5_sum <= res_5_sum + score_5_x212;
      res_6_sum <= res_6_sum + score_6_x212;
      res_7_sum <= res_7_sum + score_7_x212;
      res_8_sum <= res_8_sum + score_8_x212;
      res_9_sum <= res_9_sum + score_9_x212;
   end
   else if(res_done_x213) begin
      res_0_sum <= res_0_sum + score_0_x213;
      res_1_sum <= res_1_sum + score_1_x213;
      res_2_sum <= res_2_sum + score_2_x213;
      res_3_sum <= res_3_sum + score_3_x213;
      res_4_sum <= res_4_sum + score_4_x213;
      res_5_sum <= res_5_sum + score_5_x213;
      res_6_sum <= res_6_sum + score_6_x213;
      res_7_sum <= res_7_sum + score_7_x213;
      res_8_sum <= res_8_sum + score_8_x213;
      res_9_sum <= res_9_sum + score_9_x213;
   end
   else if(res_done_x214) begin
      res_0_sum <= res_0_sum + score_0_x214;
      res_1_sum <= res_1_sum + score_1_x214;
      res_2_sum <= res_2_sum + score_2_x214;
      res_3_sum <= res_3_sum + score_3_x214;
      res_4_sum <= res_4_sum + score_4_x214;
      res_5_sum <= res_5_sum + score_5_x214;
      res_6_sum <= res_6_sum + score_6_x214;
      res_7_sum <= res_7_sum + score_7_x214;
      res_8_sum <= res_8_sum + score_8_x214;
      res_9_sum <= res_9_sum + score_9_x214;
   end
   else if(res_done_x215) begin
      res_0_sum <= res_0_sum + score_0_x215;
      res_1_sum <= res_1_sum + score_1_x215;
      res_2_sum <= res_2_sum + score_2_x215;
      res_3_sum <= res_3_sum + score_3_x215;
      res_4_sum <= res_4_sum + score_4_x215;
      res_5_sum <= res_5_sum + score_5_x215;
      res_6_sum <= res_6_sum + score_6_x215;
      res_7_sum <= res_7_sum + score_7_x215;
      res_8_sum <= res_8_sum + score_8_x215;
      res_9_sum <= res_9_sum + score_9_x215;
   end
   else if(res_done_x216) begin
      res_0_sum <= res_0_sum + score_0_x216;
      res_1_sum <= res_1_sum + score_1_x216;
      res_2_sum <= res_2_sum + score_2_x216;
      res_3_sum <= res_3_sum + score_3_x216;
      res_4_sum <= res_4_sum + score_4_x216;
      res_5_sum <= res_5_sum + score_5_x216;
      res_6_sum <= res_6_sum + score_6_x216;
      res_7_sum <= res_7_sum + score_7_x216;
      res_8_sum <= res_8_sum + score_8_x216;
      res_9_sum <= res_9_sum + score_9_x216;
   end
   else if(res_done_x217) begin
      res_0_sum <= res_0_sum + score_0_x217;
      res_1_sum <= res_1_sum + score_1_x217;
      res_2_sum <= res_2_sum + score_2_x217;
      res_3_sum <= res_3_sum + score_3_x217;
      res_4_sum <= res_4_sum + score_4_x217;
      res_5_sum <= res_5_sum + score_5_x217;
      res_6_sum <= res_6_sum + score_6_x217;
      res_7_sum <= res_7_sum + score_7_x217;
      res_8_sum <= res_8_sum + score_8_x217;
      res_9_sum <= res_9_sum + score_9_x217;
   end
   else if(res_done_x218) begin
      res_0_sum <= res_0_sum + score_0_x218;
      res_1_sum <= res_1_sum + score_1_x218;
      res_2_sum <= res_2_sum + score_2_x218;
      res_3_sum <= res_3_sum + score_3_x218;
      res_4_sum <= res_4_sum + score_4_x218;
      res_5_sum <= res_5_sum + score_5_x218;
      res_6_sum <= res_6_sum + score_6_x218;
      res_7_sum <= res_7_sum + score_7_x218;
      res_8_sum <= res_8_sum + score_8_x218;
      res_9_sum <= res_9_sum + score_9_x218;
   end
   else if(res_done_x219) begin
      res_0_sum <= res_0_sum + score_0_x219;
      res_1_sum <= res_1_sum + score_1_x219;
      res_2_sum <= res_2_sum + score_2_x219;
      res_3_sum <= res_3_sum + score_3_x219;
      res_4_sum <= res_4_sum + score_4_x219;
      res_5_sum <= res_5_sum + score_5_x219;
      res_6_sum <= res_6_sum + score_6_x219;
      res_7_sum <= res_7_sum + score_7_x219;
      res_8_sum <= res_8_sum + score_8_x219;
      res_9_sum <= res_9_sum + score_9_x219;
   end
   else if(res_done_x220) begin
      res_0_sum <= res_0_sum + score_0_x220;
      res_1_sum <= res_1_sum + score_1_x220;
      res_2_sum <= res_2_sum + score_2_x220;
      res_3_sum <= res_3_sum + score_3_x220;
      res_4_sum <= res_4_sum + score_4_x220;
      res_5_sum <= res_5_sum + score_5_x220;
      res_6_sum <= res_6_sum + score_6_x220;
      res_7_sum <= res_7_sum + score_7_x220;
      res_8_sum <= res_8_sum + score_8_x220;
      res_9_sum <= res_9_sum + score_9_x220;
   end
   else if(res_done_x221) begin
      res_0_sum <= res_0_sum + score_0_x221;
      res_1_sum <= res_1_sum + score_1_x221;
      res_2_sum <= res_2_sum + score_2_x221;
      res_3_sum <= res_3_sum + score_3_x221;
      res_4_sum <= res_4_sum + score_4_x221;
      res_5_sum <= res_5_sum + score_5_x221;
      res_6_sum <= res_6_sum + score_6_x221;
      res_7_sum <= res_7_sum + score_7_x221;
      res_8_sum <= res_8_sum + score_8_x221;
      res_9_sum <= res_9_sum + score_9_x221;
   end
   else if(res_done_x222) begin
      res_0_sum <= res_0_sum + score_0_x222;
      res_1_sum <= res_1_sum + score_1_x222;
      res_2_sum <= res_2_sum + score_2_x222;
      res_3_sum <= res_3_sum + score_3_x222;
      res_4_sum <= res_4_sum + score_4_x222;
      res_5_sum <= res_5_sum + score_5_x222;
      res_6_sum <= res_6_sum + score_6_x222;
      res_7_sum <= res_7_sum + score_7_x222;
      res_8_sum <= res_8_sum + score_8_x222;
      res_9_sum <= res_9_sum + score_9_x222;
   end
   else if(res_done_x223) begin
      res_0_sum <= res_0_sum + score_0_x223;
      res_1_sum <= res_1_sum + score_1_x223;
      res_2_sum <= res_2_sum + score_2_x223;
      res_3_sum <= res_3_sum + score_3_x223;
      res_4_sum <= res_4_sum + score_4_x223;
      res_5_sum <= res_5_sum + score_5_x223;
      res_6_sum <= res_6_sum + score_6_x223;
      res_7_sum <= res_7_sum + score_7_x223;
      res_8_sum <= res_8_sum + score_8_x223;
      res_9_sum <= res_9_sum + score_9_x223;
   end
   else if(res_done_x224) begin
      res_0_sum <= res_0_sum + score_0_x224;
      res_1_sum <= res_1_sum + score_1_x224;
      res_2_sum <= res_2_sum + score_2_x224;
      res_3_sum <= res_3_sum + score_3_x224;
      res_4_sum <= res_4_sum + score_4_x224;
      res_5_sum <= res_5_sum + score_5_x224;
      res_6_sum <= res_6_sum + score_6_x224;
      res_7_sum <= res_7_sum + score_7_x224;
      res_8_sum <= res_8_sum + score_8_x224;
      res_9_sum <= res_9_sum + score_9_x224;
   end
   else if(res_done_x225) begin
      res_0_sum <= res_0_sum + score_0_x225;
      res_1_sum <= res_1_sum + score_1_x225;
      res_2_sum <= res_2_sum + score_2_x225;
      res_3_sum <= res_3_sum + score_3_x225;
      res_4_sum <= res_4_sum + score_4_x225;
      res_5_sum <= res_5_sum + score_5_x225;
      res_6_sum <= res_6_sum + score_6_x225;
      res_7_sum <= res_7_sum + score_7_x225;
      res_8_sum <= res_8_sum + score_8_x225;
      res_9_sum <= res_9_sum + score_9_x225;
   end
   else if(res_done_x226) begin
      res_0_sum <= res_0_sum + score_0_x226;
      res_1_sum <= res_1_sum + score_1_x226;
      res_2_sum <= res_2_sum + score_2_x226;
      res_3_sum <= res_3_sum + score_3_x226;
      res_4_sum <= res_4_sum + score_4_x226;
      res_5_sum <= res_5_sum + score_5_x226;
      res_6_sum <= res_6_sum + score_6_x226;
      res_7_sum <= res_7_sum + score_7_x226;
      res_8_sum <= res_8_sum + score_8_x226;
      res_9_sum <= res_9_sum + score_9_x226;
   end
   else if(res_done_x227) begin
      res_0_sum <= res_0_sum + score_0_x227;
      res_1_sum <= res_1_sum + score_1_x227;
      res_2_sum <= res_2_sum + score_2_x227;
      res_3_sum <= res_3_sum + score_3_x227;
      res_4_sum <= res_4_sum + score_4_x227;
      res_5_sum <= res_5_sum + score_5_x227;
      res_6_sum <= res_6_sum + score_6_x227;
      res_7_sum <= res_7_sum + score_7_x227;
      res_8_sum <= res_8_sum + score_8_x227;
      res_9_sum <= res_9_sum + score_9_x227;
   end
   else if(res_done_x228) begin
      res_0_sum <= res_0_sum + score_0_x228;
      res_1_sum <= res_1_sum + score_1_x228;
      res_2_sum <= res_2_sum + score_2_x228;
      res_3_sum <= res_3_sum + score_3_x228;
      res_4_sum <= res_4_sum + score_4_x228;
      res_5_sum <= res_5_sum + score_5_x228;
      res_6_sum <= res_6_sum + score_6_x228;
      res_7_sum <= res_7_sum + score_7_x228;
      res_8_sum <= res_8_sum + score_8_x228;
      res_9_sum <= res_9_sum + score_9_x228;
   end
   else if(res_done_x229) begin
      res_0_sum <= res_0_sum + score_0_x229;
      res_1_sum <= res_1_sum + score_1_x229;
      res_2_sum <= res_2_sum + score_2_x229;
      res_3_sum <= res_3_sum + score_3_x229;
      res_4_sum <= res_4_sum + score_4_x229;
      res_5_sum <= res_5_sum + score_5_x229;
      res_6_sum <= res_6_sum + score_6_x229;
      res_7_sum <= res_7_sum + score_7_x229;
      res_8_sum <= res_8_sum + score_8_x229;
      res_9_sum <= res_9_sum + score_9_x229;
   end
   else if(res_done_x230) begin
      res_0_sum <= res_0_sum + score_0_x230;
      res_1_sum <= res_1_sum + score_1_x230;
      res_2_sum <= res_2_sum + score_2_x230;
      res_3_sum <= res_3_sum + score_3_x230;
      res_4_sum <= res_4_sum + score_4_x230;
      res_5_sum <= res_5_sum + score_5_x230;
      res_6_sum <= res_6_sum + score_6_x230;
      res_7_sum <= res_7_sum + score_7_x230;
      res_8_sum <= res_8_sum + score_8_x230;
      res_9_sum <= res_9_sum + score_9_x230;
   end
   else if(res_done_x231) begin
      res_0_sum <= res_0_sum + score_0_x231;
      res_1_sum <= res_1_sum + score_1_x231;
      res_2_sum <= res_2_sum + score_2_x231;
      res_3_sum <= res_3_sum + score_3_x231;
      res_4_sum <= res_4_sum + score_4_x231;
      res_5_sum <= res_5_sum + score_5_x231;
      res_6_sum <= res_6_sum + score_6_x231;
      res_7_sum <= res_7_sum + score_7_x231;
      res_8_sum <= res_8_sum + score_8_x231;
      res_9_sum <= res_9_sum + score_9_x231;
   end
   else if(res_done_x232) begin
      res_0_sum <= res_0_sum + score_0_x232;
      res_1_sum <= res_1_sum + score_1_x232;
      res_2_sum <= res_2_sum + score_2_x232;
      res_3_sum <= res_3_sum + score_3_x232;
      res_4_sum <= res_4_sum + score_4_x232;
      res_5_sum <= res_5_sum + score_5_x232;
      res_6_sum <= res_6_sum + score_6_x232;
      res_7_sum <= res_7_sum + score_7_x232;
      res_8_sum <= res_8_sum + score_8_x232;
      res_9_sum <= res_9_sum + score_9_x232;
   end
   else if(res_done_x233) begin
      res_0_sum <= res_0_sum + score_0_x233;
      res_1_sum <= res_1_sum + score_1_x233;
      res_2_sum <= res_2_sum + score_2_x233;
      res_3_sum <= res_3_sum + score_3_x233;
      res_4_sum <= res_4_sum + score_4_x233;
      res_5_sum <= res_5_sum + score_5_x233;
      res_6_sum <= res_6_sum + score_6_x233;
      res_7_sum <= res_7_sum + score_7_x233;
      res_8_sum <= res_8_sum + score_8_x233;
      res_9_sum <= res_9_sum + score_9_x233;
   end
   else if(res_done_x234) begin
      res_0_sum <= res_0_sum + score_0_x234;
      res_1_sum <= res_1_sum + score_1_x234;
      res_2_sum <= res_2_sum + score_2_x234;
      res_3_sum <= res_3_sum + score_3_x234;
      res_4_sum <= res_4_sum + score_4_x234;
      res_5_sum <= res_5_sum + score_5_x234;
      res_6_sum <= res_6_sum + score_6_x234;
      res_7_sum <= res_7_sum + score_7_x234;
      res_8_sum <= res_8_sum + score_8_x234;
      res_9_sum <= res_9_sum + score_9_x234;
   end
   else if(res_done_x235) begin
      res_0_sum <= res_0_sum + score_0_x235;
      res_1_sum <= res_1_sum + score_1_x235;
      res_2_sum <= res_2_sum + score_2_x235;
      res_3_sum <= res_3_sum + score_3_x235;
      res_4_sum <= res_4_sum + score_4_x235;
      res_5_sum <= res_5_sum + score_5_x235;
      res_6_sum <= res_6_sum + score_6_x235;
      res_7_sum <= res_7_sum + score_7_x235;
      res_8_sum <= res_8_sum + score_8_x235;
      res_9_sum <= res_9_sum + score_9_x235;
   end
   else if(res_done_x236) begin
      res_0_sum <= res_0_sum + score_0_x236;
      res_1_sum <= res_1_sum + score_1_x236;
      res_2_sum <= res_2_sum + score_2_x236;
      res_3_sum <= res_3_sum + score_3_x236;
      res_4_sum <= res_4_sum + score_4_x236;
      res_5_sum <= res_5_sum + score_5_x236;
      res_6_sum <= res_6_sum + score_6_x236;
      res_7_sum <= res_7_sum + score_7_x236;
      res_8_sum <= res_8_sum + score_8_x236;
      res_9_sum <= res_9_sum + score_9_x236;
   end
   else if(res_done_x237) begin
      res_0_sum <= res_0_sum + score_0_x237;
      res_1_sum <= res_1_sum + score_1_x237;
      res_2_sum <= res_2_sum + score_2_x237;
      res_3_sum <= res_3_sum + score_3_x237;
      res_4_sum <= res_4_sum + score_4_x237;
      res_5_sum <= res_5_sum + score_5_x237;
      res_6_sum <= res_6_sum + score_6_x237;
      res_7_sum <= res_7_sum + score_7_x237;
      res_8_sum <= res_8_sum + score_8_x237;
      res_9_sum <= res_9_sum + score_9_x237;
   end
   else if(res_done_x238) begin
      res_0_sum <= res_0_sum + score_0_x238;
      res_1_sum <= res_1_sum + score_1_x238;
      res_2_sum <= res_2_sum + score_2_x238;
      res_3_sum <= res_3_sum + score_3_x238;
      res_4_sum <= res_4_sum + score_4_x238;
      res_5_sum <= res_5_sum + score_5_x238;
      res_6_sum <= res_6_sum + score_6_x238;
      res_7_sum <= res_7_sum + score_7_x238;
      res_8_sum <= res_8_sum + score_8_x238;
      res_9_sum <= res_9_sum + score_9_x238;
   end
   else if(res_done_x239) begin
      res_0_sum <= res_0_sum + score_0_x239;
      res_1_sum <= res_1_sum + score_1_x239;
      res_2_sum <= res_2_sum + score_2_x239;
      res_3_sum <= res_3_sum + score_3_x239;
      res_4_sum <= res_4_sum + score_4_x239;
      res_5_sum <= res_5_sum + score_5_x239;
      res_6_sum <= res_6_sum + score_6_x239;
      res_7_sum <= res_7_sum + score_7_x239;
      res_8_sum <= res_8_sum + score_8_x239;
      res_9_sum <= res_9_sum + score_9_x239;
   end
   else if(res_done_x240) begin
      res_0_sum <= res_0_sum + score_0_x240;
      res_1_sum <= res_1_sum + score_1_x240;
      res_2_sum <= res_2_sum + score_2_x240;
      res_3_sum <= res_3_sum + score_3_x240;
      res_4_sum <= res_4_sum + score_4_x240;
      res_5_sum <= res_5_sum + score_5_x240;
      res_6_sum <= res_6_sum + score_6_x240;
      res_7_sum <= res_7_sum + score_7_x240;
      res_8_sum <= res_8_sum + score_8_x240;
      res_9_sum <= res_9_sum + score_9_x240;
   end
   else if(res_done_x241) begin
      res_0_sum <= res_0_sum + score_0_x241;
      res_1_sum <= res_1_sum + score_1_x241;
      res_2_sum <= res_2_sum + score_2_x241;
      res_3_sum <= res_3_sum + score_3_x241;
      res_4_sum <= res_4_sum + score_4_x241;
      res_5_sum <= res_5_sum + score_5_x241;
      res_6_sum <= res_6_sum + score_6_x241;
      res_7_sum <= res_7_sum + score_7_x241;
      res_8_sum <= res_8_sum + score_8_x241;
      res_9_sum <= res_9_sum + score_9_x241;
   end
   else if(res_done_x242) begin
      res_0_sum <= res_0_sum + score_0_x242;
      res_1_sum <= res_1_sum + score_1_x242;
      res_2_sum <= res_2_sum + score_2_x242;
      res_3_sum <= res_3_sum + score_3_x242;
      res_4_sum <= res_4_sum + score_4_x242;
      res_5_sum <= res_5_sum + score_5_x242;
      res_6_sum <= res_6_sum + score_6_x242;
      res_7_sum <= res_7_sum + score_7_x242;
      res_8_sum <= res_8_sum + score_8_x242;
      res_9_sum <= res_9_sum + score_9_x242;
   end
   else if(res_done_x243) begin
      res_0_sum <= res_0_sum + score_0_x243;
      res_1_sum <= res_1_sum + score_1_x243;
      res_2_sum <= res_2_sum + score_2_x243;
      res_3_sum <= res_3_sum + score_3_x243;
      res_4_sum <= res_4_sum + score_4_x243;
      res_5_sum <= res_5_sum + score_5_x243;
      res_6_sum <= res_6_sum + score_6_x243;
      res_7_sum <= res_7_sum + score_7_x243;
      res_8_sum <= res_8_sum + score_8_x243;
      res_9_sum <= res_9_sum + score_9_x243;
   end
   else if(res_done_x244) begin
      res_0_sum <= res_0_sum + score_0_x244;
      res_1_sum <= res_1_sum + score_1_x244;
      res_2_sum <= res_2_sum + score_2_x244;
      res_3_sum <= res_3_sum + score_3_x244;
      res_4_sum <= res_4_sum + score_4_x244;
      res_5_sum <= res_5_sum + score_5_x244;
      res_6_sum <= res_6_sum + score_6_x244;
      res_7_sum <= res_7_sum + score_7_x244;
      res_8_sum <= res_8_sum + score_8_x244;
      res_9_sum <= res_9_sum + score_9_x244;
   end
   else if(res_done_x245) begin
      res_0_sum <= res_0_sum + score_0_x245;
      res_1_sum <= res_1_sum + score_1_x245;
      res_2_sum <= res_2_sum + score_2_x245;
      res_3_sum <= res_3_sum + score_3_x245;
      res_4_sum <= res_4_sum + score_4_x245;
      res_5_sum <= res_5_sum + score_5_x245;
      res_6_sum <= res_6_sum + score_6_x245;
      res_7_sum <= res_7_sum + score_7_x245;
      res_8_sum <= res_8_sum + score_8_x245;
      res_9_sum <= res_9_sum + score_9_x245;
   end
   else if(res_done_x246) begin
      res_0_sum <= res_0_sum + score_0_x246;
      res_1_sum <= res_1_sum + score_1_x246;
      res_2_sum <= res_2_sum + score_2_x246;
      res_3_sum <= res_3_sum + score_3_x246;
      res_4_sum <= res_4_sum + score_4_x246;
      res_5_sum <= res_5_sum + score_5_x246;
      res_6_sum <= res_6_sum + score_6_x246;
      res_7_sum <= res_7_sum + score_7_x246;
      res_8_sum <= res_8_sum + score_8_x246;
      res_9_sum <= res_9_sum + score_9_x246;
   end
   else if(res_done_x247) begin
      res_0_sum <= res_0_sum + score_0_x247;
      res_1_sum <= res_1_sum + score_1_x247;
      res_2_sum <= res_2_sum + score_2_x247;
      res_3_sum <= res_3_sum + score_3_x247;
      res_4_sum <= res_4_sum + score_4_x247;
      res_5_sum <= res_5_sum + score_5_x247;
      res_6_sum <= res_6_sum + score_6_x247;
      res_7_sum <= res_7_sum + score_7_x247;
      res_8_sum <= res_8_sum + score_8_x247;
      res_9_sum <= res_9_sum + score_9_x247;
   end
   else if(res_done_x248) begin
      res_0_sum <= res_0_sum + score_0_x248;
      res_1_sum <= res_1_sum + score_1_x248;
      res_2_sum <= res_2_sum + score_2_x248;
      res_3_sum <= res_3_sum + score_3_x248;
      res_4_sum <= res_4_sum + score_4_x248;
      res_5_sum <= res_5_sum + score_5_x248;
      res_6_sum <= res_6_sum + score_6_x248;
      res_7_sum <= res_7_sum + score_7_x248;
      res_8_sum <= res_8_sum + score_8_x248;
      res_9_sum <= res_9_sum + score_9_x248;
   end
   else if(res_done_x249) begin
      res_0_sum <= res_0_sum + score_0_x249;
      res_1_sum <= res_1_sum + score_1_x249;
      res_2_sum <= res_2_sum + score_2_x249;
      res_3_sum <= res_3_sum + score_3_x249;
      res_4_sum <= res_4_sum + score_4_x249;
      res_5_sum <= res_5_sum + score_5_x249;
      res_6_sum <= res_6_sum + score_6_x249;
      res_7_sum <= res_7_sum + score_7_x249;
      res_8_sum <= res_8_sum + score_8_x249;
      res_9_sum <= res_9_sum + score_9_x249;
   end
   else if(res_done_x250) begin
      res_0_sum <= res_0_sum + score_0_x250;
      res_1_sum <= res_1_sum + score_1_x250;
      res_2_sum <= res_2_sum + score_2_x250;
      res_3_sum <= res_3_sum + score_3_x250;
      res_4_sum <= res_4_sum + score_4_x250;
      res_5_sum <= res_5_sum + score_5_x250;
      res_6_sum <= res_6_sum + score_6_x250;
      res_7_sum <= res_7_sum + score_7_x250;
      res_8_sum <= res_8_sum + score_8_x250;
      res_9_sum <= res_9_sum + score_9_x250;
   end
   else if(res_done_x251) begin
      res_0_sum <= res_0_sum + score_0_x251;
      res_1_sum <= res_1_sum + score_1_x251;
      res_2_sum <= res_2_sum + score_2_x251;
      res_3_sum <= res_3_sum + score_3_x251;
      res_4_sum <= res_4_sum + score_4_x251;
      res_5_sum <= res_5_sum + score_5_x251;
      res_6_sum <= res_6_sum + score_6_x251;
      res_7_sum <= res_7_sum + score_7_x251;
      res_8_sum <= res_8_sum + score_8_x251;
      res_9_sum <= res_9_sum + score_9_x251;
   end
   else if(res_done_x252) begin
      res_0_sum <= res_0_sum + score_0_x252;
      res_1_sum <= res_1_sum + score_1_x252;
      res_2_sum <= res_2_sum + score_2_x252;
      res_3_sum <= res_3_sum + score_3_x252;
      res_4_sum <= res_4_sum + score_4_x252;
      res_5_sum <= res_5_sum + score_5_x252;
      res_6_sum <= res_6_sum + score_6_x252;
      res_7_sum <= res_7_sum + score_7_x252;
      res_8_sum <= res_8_sum + score_8_x252;
      res_9_sum <= res_9_sum + score_9_x252;
   end
   else if(res_done_x253) begin
      res_0_sum <= res_0_sum + score_0_x253;
      res_1_sum <= res_1_sum + score_1_x253;
      res_2_sum <= res_2_sum + score_2_x253;
      res_3_sum <= res_3_sum + score_3_x253;
      res_4_sum <= res_4_sum + score_4_x253;
      res_5_sum <= res_5_sum + score_5_x253;
      res_6_sum <= res_6_sum + score_6_x253;
      res_7_sum <= res_7_sum + score_7_x253;
      res_8_sum <= res_8_sum + score_8_x253;
      res_9_sum <= res_9_sum + score_9_x253;
   end
   else if(res_done_x254) begin
      res_0_sum <= res_0_sum + score_0_x254;
      res_1_sum <= res_1_sum + score_1_x254;
      res_2_sum <= res_2_sum + score_2_x254;
      res_3_sum <= res_3_sum + score_3_x254;
      res_4_sum <= res_4_sum + score_4_x254;
      res_5_sum <= res_5_sum + score_5_x254;
      res_6_sum <= res_6_sum + score_6_x254;
      res_7_sum <= res_7_sum + score_7_x254;
      res_8_sum <= res_8_sum + score_8_x254;
      res_9_sum <= res_9_sum + score_9_x254;
   end
   else if(res_done_x255) begin
      res_0_sum <= res_0_sum + score_0_x255;
      res_1_sum <= res_1_sum + score_1_x255;
      res_2_sum <= res_2_sum + score_2_x255;
      res_3_sum <= res_3_sum + score_3_x255;
      res_4_sum <= res_4_sum + score_4_x255;
      res_5_sum <= res_5_sum + score_5_x255;
      res_6_sum <= res_6_sum + score_6_x255;
      res_7_sum <= res_7_sum + score_7_x255;
      res_8_sum <= res_8_sum + score_8_x255;
      res_9_sum <= res_9_sum + score_9_x255;
   end
   else if(res_done_x256) begin
      res_0_sum <= res_0_sum + score_0_x256;
      res_1_sum <= res_1_sum + score_1_x256;
      res_2_sum <= res_2_sum + score_2_x256;
      res_3_sum <= res_3_sum + score_3_x256;
      res_4_sum <= res_4_sum + score_4_x256;
      res_5_sum <= res_5_sum + score_5_x256;
      res_6_sum <= res_6_sum + score_6_x256;
      res_7_sum <= res_7_sum + score_7_x256;
      res_8_sum <= res_8_sum + score_8_x256;
      res_9_sum <= res_9_sum + score_9_x256;
   end
   else if(res_done_x257) begin
      res_0_sum <= res_0_sum + score_0_x257;
      res_1_sum <= res_1_sum + score_1_x257;
      res_2_sum <= res_2_sum + score_2_x257;
      res_3_sum <= res_3_sum + score_3_x257;
      res_4_sum <= res_4_sum + score_4_x257;
      res_5_sum <= res_5_sum + score_5_x257;
      res_6_sum <= res_6_sum + score_6_x257;
      res_7_sum <= res_7_sum + score_7_x257;
      res_8_sum <= res_8_sum + score_8_x257;
      res_9_sum <= res_9_sum + score_9_x257;
   end
   else if(res_done_x258) begin
      res_0_sum <= res_0_sum + score_0_x258;
      res_1_sum <= res_1_sum + score_1_x258;
      res_2_sum <= res_2_sum + score_2_x258;
      res_3_sum <= res_3_sum + score_3_x258;
      res_4_sum <= res_4_sum + score_4_x258;
      res_5_sum <= res_5_sum + score_5_x258;
      res_6_sum <= res_6_sum + score_6_x258;
      res_7_sum <= res_7_sum + score_7_x258;
      res_8_sum <= res_8_sum + score_8_x258;
      res_9_sum <= res_9_sum + score_9_x258;
   end
   else if(res_done_x259) begin
      res_0_sum <= res_0_sum + score_0_x259;
      res_1_sum <= res_1_sum + score_1_x259;
      res_2_sum <= res_2_sum + score_2_x259;
      res_3_sum <= res_3_sum + score_3_x259;
      res_4_sum <= res_4_sum + score_4_x259;
      res_5_sum <= res_5_sum + score_5_x259;
      res_6_sum <= res_6_sum + score_6_x259;
      res_7_sum <= res_7_sum + score_7_x259;
      res_8_sum <= res_8_sum + score_8_x259;
      res_9_sum <= res_9_sum + score_9_x259;
   end
   else if(res_done_x260) begin
      res_0_sum <= res_0_sum + score_0_x260;
      res_1_sum <= res_1_sum + score_1_x260;
      res_2_sum <= res_2_sum + score_2_x260;
      res_3_sum <= res_3_sum + score_3_x260;
      res_4_sum <= res_4_sum + score_4_x260;
      res_5_sum <= res_5_sum + score_5_x260;
      res_6_sum <= res_6_sum + score_6_x260;
      res_7_sum <= res_7_sum + score_7_x260;
      res_8_sum <= res_8_sum + score_8_x260;
      res_9_sum <= res_9_sum + score_9_x260;
   end
   else if(res_done_x261) begin
      res_0_sum <= res_0_sum + score_0_x261;
      res_1_sum <= res_1_sum + score_1_x261;
      res_2_sum <= res_2_sum + score_2_x261;
      res_3_sum <= res_3_sum + score_3_x261;
      res_4_sum <= res_4_sum + score_4_x261;
      res_5_sum <= res_5_sum + score_5_x261;
      res_6_sum <= res_6_sum + score_6_x261;
      res_7_sum <= res_7_sum + score_7_x261;
      res_8_sum <= res_8_sum + score_8_x261;
      res_9_sum <= res_9_sum + score_9_x261;
   end
   else if(res_done_x262) begin
      res_0_sum <= res_0_sum + score_0_x262;
      res_1_sum <= res_1_sum + score_1_x262;
      res_2_sum <= res_2_sum + score_2_x262;
      res_3_sum <= res_3_sum + score_3_x262;
      res_4_sum <= res_4_sum + score_4_x262;
      res_5_sum <= res_5_sum + score_5_x262;
      res_6_sum <= res_6_sum + score_6_x262;
      res_7_sum <= res_7_sum + score_7_x262;
      res_8_sum <= res_8_sum + score_8_x262;
      res_9_sum <= res_9_sum + score_9_x262;
   end
   else if(res_done_x263) begin
      res_0_sum <= res_0_sum + score_0_x263;
      res_1_sum <= res_1_sum + score_1_x263;
      res_2_sum <= res_2_sum + score_2_x263;
      res_3_sum <= res_3_sum + score_3_x263;
      res_4_sum <= res_4_sum + score_4_x263;
      res_5_sum <= res_5_sum + score_5_x263;
      res_6_sum <= res_6_sum + score_6_x263;
      res_7_sum <= res_7_sum + score_7_x263;
      res_8_sum <= res_8_sum + score_8_x263;
      res_9_sum <= res_9_sum + score_9_x263;
   end
   else if(res_done_x264) begin
      res_0_sum <= res_0_sum + score_0_x264;
      res_1_sum <= res_1_sum + score_1_x264;
      res_2_sum <= res_2_sum + score_2_x264;
      res_3_sum <= res_3_sum + score_3_x264;
      res_4_sum <= res_4_sum + score_4_x264;
      res_5_sum <= res_5_sum + score_5_x264;
      res_6_sum <= res_6_sum + score_6_x264;
      res_7_sum <= res_7_sum + score_7_x264;
      res_8_sum <= res_8_sum + score_8_x264;
      res_9_sum <= res_9_sum + score_9_x264;
   end
   else if(res_done_x265) begin
      res_0_sum <= res_0_sum + score_0_x265;
      res_1_sum <= res_1_sum + score_1_x265;
      res_2_sum <= res_2_sum + score_2_x265;
      res_3_sum <= res_3_sum + score_3_x265;
      res_4_sum <= res_4_sum + score_4_x265;
      res_5_sum <= res_5_sum + score_5_x265;
      res_6_sum <= res_6_sum + score_6_x265;
      res_7_sum <= res_7_sum + score_7_x265;
      res_8_sum <= res_8_sum + score_8_x265;
      res_9_sum <= res_9_sum + score_9_x265;
   end
   else if(res_done_x266) begin
      res_0_sum <= res_0_sum + score_0_x266;
      res_1_sum <= res_1_sum + score_1_x266;
      res_2_sum <= res_2_sum + score_2_x266;
      res_3_sum <= res_3_sum + score_3_x266;
      res_4_sum <= res_4_sum + score_4_x266;
      res_5_sum <= res_5_sum + score_5_x266;
      res_6_sum <= res_6_sum + score_6_x266;
      res_7_sum <= res_7_sum + score_7_x266;
      res_8_sum <= res_8_sum + score_8_x266;
      res_9_sum <= res_9_sum + score_9_x266;
   end
   else if(res_done_x267) begin
      res_0_sum <= res_0_sum + score_0_x267;
      res_1_sum <= res_1_sum + score_1_x267;
      res_2_sum <= res_2_sum + score_2_x267;
      res_3_sum <= res_3_sum + score_3_x267;
      res_4_sum <= res_4_sum + score_4_x267;
      res_5_sum <= res_5_sum + score_5_x267;
      res_6_sum <= res_6_sum + score_6_x267;
      res_7_sum <= res_7_sum + score_7_x267;
      res_8_sum <= res_8_sum + score_8_x267;
      res_9_sum <= res_9_sum + score_9_x267;
   end
   else if(res_done_x268) begin
      res_0_sum <= res_0_sum + score_0_x268;
      res_1_sum <= res_1_sum + score_1_x268;
      res_2_sum <= res_2_sum + score_2_x268;
      res_3_sum <= res_3_sum + score_3_x268;
      res_4_sum <= res_4_sum + score_4_x268;
      res_5_sum <= res_5_sum + score_5_x268;
      res_6_sum <= res_6_sum + score_6_x268;
      res_7_sum <= res_7_sum + score_7_x268;
      res_8_sum <= res_8_sum + score_8_x268;
      res_9_sum <= res_9_sum + score_9_x268;
   end
   else if(res_done_x269) begin
      res_0_sum <= res_0_sum + score_0_x269;
      res_1_sum <= res_1_sum + score_1_x269;
      res_2_sum <= res_2_sum + score_2_x269;
      res_3_sum <= res_3_sum + score_3_x269;
      res_4_sum <= res_4_sum + score_4_x269;
      res_5_sum <= res_5_sum + score_5_x269;
      res_6_sum <= res_6_sum + score_6_x269;
      res_7_sum <= res_7_sum + score_7_x269;
      res_8_sum <= res_8_sum + score_8_x269;
      res_9_sum <= res_9_sum + score_9_x269;
   end
   else if(res_done_x270) begin
      res_0_sum <= res_0_sum + score_0_x270;
      res_1_sum <= res_1_sum + score_1_x270;
      res_2_sum <= res_2_sum + score_2_x270;
      res_3_sum <= res_3_sum + score_3_x270;
      res_4_sum <= res_4_sum + score_4_x270;
      res_5_sum <= res_5_sum + score_5_x270;
      res_6_sum <= res_6_sum + score_6_x270;
      res_7_sum <= res_7_sum + score_7_x270;
      res_8_sum <= res_8_sum + score_8_x270;
      res_9_sum <= res_9_sum + score_9_x270;
   end
   else if(res_done_x271) begin
      res_0_sum <= res_0_sum + score_0_x271;
      res_1_sum <= res_1_sum + score_1_x271;
      res_2_sum <= res_2_sum + score_2_x271;
      res_3_sum <= res_3_sum + score_3_x271;
      res_4_sum <= res_4_sum + score_4_x271;
      res_5_sum <= res_5_sum + score_5_x271;
      res_6_sum <= res_6_sum + score_6_x271;
      res_7_sum <= res_7_sum + score_7_x271;
      res_8_sum <= res_8_sum + score_8_x271;
      res_9_sum <= res_9_sum + score_9_x271;
   end
   else if(res_done_x272) begin
      res_0_sum <= res_0_sum + score_0_x272;
      res_1_sum <= res_1_sum + score_1_x272;
      res_2_sum <= res_2_sum + score_2_x272;
      res_3_sum <= res_3_sum + score_3_x272;
      res_4_sum <= res_4_sum + score_4_x272;
      res_5_sum <= res_5_sum + score_5_x272;
      res_6_sum <= res_6_sum + score_6_x272;
      res_7_sum <= res_7_sum + score_7_x272;
      res_8_sum <= res_8_sum + score_8_x272;
      res_9_sum <= res_9_sum + score_9_x272;
   end
   else if(res_done_x273) begin
      res_0_sum <= res_0_sum + score_0_x273;
      res_1_sum <= res_1_sum + score_1_x273;
      res_2_sum <= res_2_sum + score_2_x273;
      res_3_sum <= res_3_sum + score_3_x273;
      res_4_sum <= res_4_sum + score_4_x273;
      res_5_sum <= res_5_sum + score_5_x273;
      res_6_sum <= res_6_sum + score_6_x273;
      res_7_sum <= res_7_sum + score_7_x273;
      res_8_sum <= res_8_sum + score_8_x273;
      res_9_sum <= res_9_sum + score_9_x273;
   end
   else if(res_done_x274) begin
      res_0_sum <= res_0_sum + score_0_x274;
      res_1_sum <= res_1_sum + score_1_x274;
      res_2_sum <= res_2_sum + score_2_x274;
      res_3_sum <= res_3_sum + score_3_x274;
      res_4_sum <= res_4_sum + score_4_x274;
      res_5_sum <= res_5_sum + score_5_x274;
      res_6_sum <= res_6_sum + score_6_x274;
      res_7_sum <= res_7_sum + score_7_x274;
      res_8_sum <= res_8_sum + score_8_x274;
      res_9_sum <= res_9_sum + score_9_x274;
   end
   else if(res_done_x275) begin
      res_0_sum <= res_0_sum + score_0_x275;
      res_1_sum <= res_1_sum + score_1_x275;
      res_2_sum <= res_2_sum + score_2_x275;
      res_3_sum <= res_3_sum + score_3_x275;
      res_4_sum <= res_4_sum + score_4_x275;
      res_5_sum <= res_5_sum + score_5_x275;
      res_6_sum <= res_6_sum + score_6_x275;
      res_7_sum <= res_7_sum + score_7_x275;
      res_8_sum <= res_8_sum + score_8_x275;
      res_9_sum <= res_9_sum + score_9_x275;
   end
   else if(res_done_x276) begin
      res_0_sum <= res_0_sum + score_0_x276;
      res_1_sum <= res_1_sum + score_1_x276;
      res_2_sum <= res_2_sum + score_2_x276;
      res_3_sum <= res_3_sum + score_3_x276;
      res_4_sum <= res_4_sum + score_4_x276;
      res_5_sum <= res_5_sum + score_5_x276;
      res_6_sum <= res_6_sum + score_6_x276;
      res_7_sum <= res_7_sum + score_7_x276;
      res_8_sum <= res_8_sum + score_8_x276;
      res_9_sum <= res_9_sum + score_9_x276;
   end
   else if(res_done_x277) begin
      res_0_sum <= res_0_sum + score_0_x277;
      res_1_sum <= res_1_sum + score_1_x277;
      res_2_sum <= res_2_sum + score_2_x277;
      res_3_sum <= res_3_sum + score_3_x277;
      res_4_sum <= res_4_sum + score_4_x277;
      res_5_sum <= res_5_sum + score_5_x277;
      res_6_sum <= res_6_sum + score_6_x277;
      res_7_sum <= res_7_sum + score_7_x277;
      res_8_sum <= res_8_sum + score_8_x277;
      res_9_sum <= res_9_sum + score_9_x277;
   end
   else if(res_done_x278) begin
      res_0_sum <= res_0_sum + score_0_x278;
      res_1_sum <= res_1_sum + score_1_x278;
      res_2_sum <= res_2_sum + score_2_x278;
      res_3_sum <= res_3_sum + score_3_x278;
      res_4_sum <= res_4_sum + score_4_x278;
      res_5_sum <= res_5_sum + score_5_x278;
      res_6_sum <= res_6_sum + score_6_x278;
      res_7_sum <= res_7_sum + score_7_x278;
      res_8_sum <= res_8_sum + score_8_x278;
      res_9_sum <= res_9_sum + score_9_x278;
   end
   else if(res_done_x279) begin
      res_0_sum <= res_0_sum + score_0_x279;
      res_1_sum <= res_1_sum + score_1_x279;
      res_2_sum <= res_2_sum + score_2_x279;
      res_3_sum <= res_3_sum + score_3_x279;
      res_4_sum <= res_4_sum + score_4_x279;
      res_5_sum <= res_5_sum + score_5_x279;
      res_6_sum <= res_6_sum + score_6_x279;
      res_7_sum <= res_7_sum + score_7_x279;
      res_8_sum <= res_8_sum + score_8_x279;
      res_9_sum <= res_9_sum + score_9_x279;
   end
   else if(res_done_x280) begin
      res_0_sum <= res_0_sum + score_0_x280;
      res_1_sum <= res_1_sum + score_1_x280;
      res_2_sum <= res_2_sum + score_2_x280;
      res_3_sum <= res_3_sum + score_3_x280;
      res_4_sum <= res_4_sum + score_4_x280;
      res_5_sum <= res_5_sum + score_5_x280;
      res_6_sum <= res_6_sum + score_6_x280;
      res_7_sum <= res_7_sum + score_7_x280;
      res_8_sum <= res_8_sum + score_8_x280;
      res_9_sum <= res_9_sum + score_9_x280;
   end
   else if(res_done_x281) begin
      res_0_sum <= res_0_sum + score_0_x281;
      res_1_sum <= res_1_sum + score_1_x281;
      res_2_sum <= res_2_sum + score_2_x281;
      res_3_sum <= res_3_sum + score_3_x281;
      res_4_sum <= res_4_sum + score_4_x281;
      res_5_sum <= res_5_sum + score_5_x281;
      res_6_sum <= res_6_sum + score_6_x281;
      res_7_sum <= res_7_sum + score_7_x281;
      res_8_sum <= res_8_sum + score_8_x281;
      res_9_sum <= res_9_sum + score_9_x281;
   end
   else if(res_done_x282) begin
      res_0_sum <= res_0_sum + score_0_x282;
      res_1_sum <= res_1_sum + score_1_x282;
      res_2_sum <= res_2_sum + score_2_x282;
      res_3_sum <= res_3_sum + score_3_x282;
      res_4_sum <= res_4_sum + score_4_x282;
      res_5_sum <= res_5_sum + score_5_x282;
      res_6_sum <= res_6_sum + score_6_x282;
      res_7_sum <= res_7_sum + score_7_x282;
      res_8_sum <= res_8_sum + score_8_x282;
      res_9_sum <= res_9_sum + score_9_x282;
   end
   else if(res_done_x283) begin
      res_0_sum <= res_0_sum + score_0_x283;
      res_1_sum <= res_1_sum + score_1_x283;
      res_2_sum <= res_2_sum + score_2_x283;
      res_3_sum <= res_3_sum + score_3_x283;
      res_4_sum <= res_4_sum + score_4_x283;
      res_5_sum <= res_5_sum + score_5_x283;
      res_6_sum <= res_6_sum + score_6_x283;
      res_7_sum <= res_7_sum + score_7_x283;
      res_8_sum <= res_8_sum + score_8_x283;
      res_9_sum <= res_9_sum + score_9_x283;
   end
   else if(res_done_x284) begin
      res_0_sum <= res_0_sum + score_0_x284;
      res_1_sum <= res_1_sum + score_1_x284;
      res_2_sum <= res_2_sum + score_2_x284;
      res_3_sum <= res_3_sum + score_3_x284;
      res_4_sum <= res_4_sum + score_4_x284;
      res_5_sum <= res_5_sum + score_5_x284;
      res_6_sum <= res_6_sum + score_6_x284;
      res_7_sum <= res_7_sum + score_7_x284;
      res_8_sum <= res_8_sum + score_8_x284;
      res_9_sum <= res_9_sum + score_9_x284;
   end
   else if(res_done_x285) begin
      res_0_sum <= res_0_sum + score_0_x285;
      res_1_sum <= res_1_sum + score_1_x285;
      res_2_sum <= res_2_sum + score_2_x285;
      res_3_sum <= res_3_sum + score_3_x285;
      res_4_sum <= res_4_sum + score_4_x285;
      res_5_sum <= res_5_sum + score_5_x285;
      res_6_sum <= res_6_sum + score_6_x285;
      res_7_sum <= res_7_sum + score_7_x285;
      res_8_sum <= res_8_sum + score_8_x285;
      res_9_sum <= res_9_sum + score_9_x285;
   end
   else if(res_done_x286) begin
      res_0_sum <= res_0_sum + score_0_x286;
      res_1_sum <= res_1_sum + score_1_x286;
      res_2_sum <= res_2_sum + score_2_x286;
      res_3_sum <= res_3_sum + score_3_x286;
      res_4_sum <= res_4_sum + score_4_x286;
      res_5_sum <= res_5_sum + score_5_x286;
      res_6_sum <= res_6_sum + score_6_x286;
      res_7_sum <= res_7_sum + score_7_x286;
      res_8_sum <= res_8_sum + score_8_x286;
      res_9_sum <= res_9_sum + score_9_x286;
   end
   else if(res_done_x287) begin
      res_0_sum <= res_0_sum + score_0_x287;
      res_1_sum <= res_1_sum + score_1_x287;
      res_2_sum <= res_2_sum + score_2_x287;
      res_3_sum <= res_3_sum + score_3_x287;
      res_4_sum <= res_4_sum + score_4_x287;
      res_5_sum <= res_5_sum + score_5_x287;
      res_6_sum <= res_6_sum + score_6_x287;
      res_7_sum <= res_7_sum + score_7_x287;
      res_8_sum <= res_8_sum + score_8_x287;
      res_9_sum <= res_9_sum + score_9_x287;
   end
   else if(res_done_x288) begin
      res_0_sum <= res_0_sum + score_0_x288;
      res_1_sum <= res_1_sum + score_1_x288;
      res_2_sum <= res_2_sum + score_2_x288;
      res_3_sum <= res_3_sum + score_3_x288;
      res_4_sum <= res_4_sum + score_4_x288;
      res_5_sum <= res_5_sum + score_5_x288;
      res_6_sum <= res_6_sum + score_6_x288;
      res_7_sum <= res_7_sum + score_7_x288;
      res_8_sum <= res_8_sum + score_8_x288;
      res_9_sum <= res_9_sum + score_9_x288;
   end
   else if(res_done_x289) begin
      res_0_sum <= res_0_sum + score_0_x289;
      res_1_sum <= res_1_sum + score_1_x289;
      res_2_sum <= res_2_sum + score_2_x289;
      res_3_sum <= res_3_sum + score_3_x289;
      res_4_sum <= res_4_sum + score_4_x289;
      res_5_sum <= res_5_sum + score_5_x289;
      res_6_sum <= res_6_sum + score_6_x289;
      res_7_sum <= res_7_sum + score_7_x289;
      res_8_sum <= res_8_sum + score_8_x289;
      res_9_sum <= res_9_sum + score_9_x289;
   end
   else if(res_done_x290) begin
      res_0_sum <= res_0_sum + score_0_x290;
      res_1_sum <= res_1_sum + score_1_x290;
      res_2_sum <= res_2_sum + score_2_x290;
      res_3_sum <= res_3_sum + score_3_x290;
      res_4_sum <= res_4_sum + score_4_x290;
      res_5_sum <= res_5_sum + score_5_x290;
      res_6_sum <= res_6_sum + score_6_x290;
      res_7_sum <= res_7_sum + score_7_x290;
      res_8_sum <= res_8_sum + score_8_x290;
      res_9_sum <= res_9_sum + score_9_x290;
   end
   else if(res_done_x291) begin
      res_0_sum <= res_0_sum + score_0_x291;
      res_1_sum <= res_1_sum + score_1_x291;
      res_2_sum <= res_2_sum + score_2_x291;
      res_3_sum <= res_3_sum + score_3_x291;
      res_4_sum <= res_4_sum + score_4_x291;
      res_5_sum <= res_5_sum + score_5_x291;
      res_6_sum <= res_6_sum + score_6_x291;
      res_7_sum <= res_7_sum + score_7_x291;
      res_8_sum <= res_8_sum + score_8_x291;
      res_9_sum <= res_9_sum + score_9_x291;
   end
   else if(res_done_x292) begin
      res_0_sum <= res_0_sum + score_0_x292;
      res_1_sum <= res_1_sum + score_1_x292;
      res_2_sum <= res_2_sum + score_2_x292;
      res_3_sum <= res_3_sum + score_3_x292;
      res_4_sum <= res_4_sum + score_4_x292;
      res_5_sum <= res_5_sum + score_5_x292;
      res_6_sum <= res_6_sum + score_6_x292;
      res_7_sum <= res_7_sum + score_7_x292;
      res_8_sum <= res_8_sum + score_8_x292;
      res_9_sum <= res_9_sum + score_9_x292;
   end
   else if(res_done_x293) begin
      res_0_sum <= res_0_sum + score_0_x293;
      res_1_sum <= res_1_sum + score_1_x293;
      res_2_sum <= res_2_sum + score_2_x293;
      res_3_sum <= res_3_sum + score_3_x293;
      res_4_sum <= res_4_sum + score_4_x293;
      res_5_sum <= res_5_sum + score_5_x293;
      res_6_sum <= res_6_sum + score_6_x293;
      res_7_sum <= res_7_sum + score_7_x293;
      res_8_sum <= res_8_sum + score_8_x293;
      res_9_sum <= res_9_sum + score_9_x293;
   end
   else if(res_done_x294) begin
      res_0_sum <= res_0_sum + score_0_x294;
      res_1_sum <= res_1_sum + score_1_x294;
      res_2_sum <= res_2_sum + score_2_x294;
      res_3_sum <= res_3_sum + score_3_x294;
      res_4_sum <= res_4_sum + score_4_x294;
      res_5_sum <= res_5_sum + score_5_x294;
      res_6_sum <= res_6_sum + score_6_x294;
      res_7_sum <= res_7_sum + score_7_x294;
      res_8_sum <= res_8_sum + score_8_x294;
      res_9_sum <= res_9_sum + score_9_x294;
   end
   else if(res_done_x295) begin
      res_0_sum <= res_0_sum + score_0_x295;
      res_1_sum <= res_1_sum + score_1_x295;
      res_2_sum <= res_2_sum + score_2_x295;
      res_3_sum <= res_3_sum + score_3_x295;
      res_4_sum <= res_4_sum + score_4_x295;
      res_5_sum <= res_5_sum + score_5_x295;
      res_6_sum <= res_6_sum + score_6_x295;
      res_7_sum <= res_7_sum + score_7_x295;
      res_8_sum <= res_8_sum + score_8_x295;
      res_9_sum <= res_9_sum + score_9_x295;
   end
   else if(res_done_x296) begin
      res_0_sum <= res_0_sum + score_0_x296;
      res_1_sum <= res_1_sum + score_1_x296;
      res_2_sum <= res_2_sum + score_2_x296;
      res_3_sum <= res_3_sum + score_3_x296;
      res_4_sum <= res_4_sum + score_4_x296;
      res_5_sum <= res_5_sum + score_5_x296;
      res_6_sum <= res_6_sum + score_6_x296;
      res_7_sum <= res_7_sum + score_7_x296;
      res_8_sum <= res_8_sum + score_8_x296;
      res_9_sum <= res_9_sum + score_9_x296;
   end
   else if(res_done_x297) begin
      res_0_sum <= res_0_sum + score_0_x297;
      res_1_sum <= res_1_sum + score_1_x297;
      res_2_sum <= res_2_sum + score_2_x297;
      res_3_sum <= res_3_sum + score_3_x297;
      res_4_sum <= res_4_sum + score_4_x297;
      res_5_sum <= res_5_sum + score_5_x297;
      res_6_sum <= res_6_sum + score_6_x297;
      res_7_sum <= res_7_sum + score_7_x297;
      res_8_sum <= res_8_sum + score_8_x297;
      res_9_sum <= res_9_sum + score_9_x297;
   end
   else if(res_done_x298) begin
      res_0_sum <= res_0_sum + score_0_x298;
      res_1_sum <= res_1_sum + score_1_x298;
      res_2_sum <= res_2_sum + score_2_x298;
      res_3_sum <= res_3_sum + score_3_x298;
      res_4_sum <= res_4_sum + score_4_x298;
      res_5_sum <= res_5_sum + score_5_x298;
      res_6_sum <= res_6_sum + score_6_x298;
      res_7_sum <= res_7_sum + score_7_x298;
      res_8_sum <= res_8_sum + score_8_x298;
      res_9_sum <= res_9_sum + score_9_x298;
   end
   else if(res_done_x299) begin
      res_0_sum <= res_0_sum + score_0_x299;
      res_1_sum <= res_1_sum + score_1_x299;
      res_2_sum <= res_2_sum + score_2_x299;
      res_3_sum <= res_3_sum + score_3_x299;
      res_4_sum <= res_4_sum + score_4_x299;
      res_5_sum <= res_5_sum + score_5_x299;
      res_6_sum <= res_6_sum + score_6_x299;
      res_7_sum <= res_7_sum + score_7_x299;
      res_8_sum <= res_8_sum + score_8_x299;
      res_9_sum <= res_9_sum + score_9_x299;
   end
   else if(res_done_x300) begin
      res_0_sum <= res_0_sum + score_0_x300;
      res_1_sum <= res_1_sum + score_1_x300;
      res_2_sum <= res_2_sum + score_2_x300;
      res_3_sum <= res_3_sum + score_3_x300;
      res_4_sum <= res_4_sum + score_4_x300;
      res_5_sum <= res_5_sum + score_5_x300;
      res_6_sum <= res_6_sum + score_6_x300;
      res_7_sum <= res_7_sum + score_7_x300;
      res_8_sum <= res_8_sum + score_8_x300;
      res_9_sum <= res_9_sum + score_9_x300;
   end
   else if(res_done_x301) begin
      res_0_sum <= res_0_sum + score_0_x301;
      res_1_sum <= res_1_sum + score_1_x301;
      res_2_sum <= res_2_sum + score_2_x301;
      res_3_sum <= res_3_sum + score_3_x301;
      res_4_sum <= res_4_sum + score_4_x301;
      res_5_sum <= res_5_sum + score_5_x301;
      res_6_sum <= res_6_sum + score_6_x301;
      res_7_sum <= res_7_sum + score_7_x301;
      res_8_sum <= res_8_sum + score_8_x301;
      res_9_sum <= res_9_sum + score_9_x301;
   end
   else if(res_done_x302) begin
      res_0_sum <= res_0_sum + score_0_x302;
      res_1_sum <= res_1_sum + score_1_x302;
      res_2_sum <= res_2_sum + score_2_x302;
      res_3_sum <= res_3_sum + score_3_x302;
      res_4_sum <= res_4_sum + score_4_x302;
      res_5_sum <= res_5_sum + score_5_x302;
      res_6_sum <= res_6_sum + score_6_x302;
      res_7_sum <= res_7_sum + score_7_x302;
      res_8_sum <= res_8_sum + score_8_x302;
      res_9_sum <= res_9_sum + score_9_x302;
   end
   else if(res_done_x303) begin
      res_0_sum <= res_0_sum + score_0_x303;
      res_1_sum <= res_1_sum + score_1_x303;
      res_2_sum <= res_2_sum + score_2_x303;
      res_3_sum <= res_3_sum + score_3_x303;
      res_4_sum <= res_4_sum + score_4_x303;
      res_5_sum <= res_5_sum + score_5_x303;
      res_6_sum <= res_6_sum + score_6_x303;
      res_7_sum <= res_7_sum + score_7_x303;
      res_8_sum <= res_8_sum + score_8_x303;
      res_9_sum <= res_9_sum + score_9_x303;
   end
   else if(res_done_x304) begin
      res_0_sum <= res_0_sum + score_0_x304;
      res_1_sum <= res_1_sum + score_1_x304;
      res_2_sum <= res_2_sum + score_2_x304;
      res_3_sum <= res_3_sum + score_3_x304;
      res_4_sum <= res_4_sum + score_4_x304;
      res_5_sum <= res_5_sum + score_5_x304;
      res_6_sum <= res_6_sum + score_6_x304;
      res_7_sum <= res_7_sum + score_7_x304;
      res_8_sum <= res_8_sum + score_8_x304;
      res_9_sum <= res_9_sum + score_9_x304;
   end
   else if(res_done_x305) begin
      res_0_sum <= res_0_sum + score_0_x305;
      res_1_sum <= res_1_sum + score_1_x305;
      res_2_sum <= res_2_sum + score_2_x305;
      res_3_sum <= res_3_sum + score_3_x305;
      res_4_sum <= res_4_sum + score_4_x305;
      res_5_sum <= res_5_sum + score_5_x305;
      res_6_sum <= res_6_sum + score_6_x305;
      res_7_sum <= res_7_sum + score_7_x305;
      res_8_sum <= res_8_sum + score_8_x305;
      res_9_sum <= res_9_sum + score_9_x305;
   end
   else if(res_done_x306) begin
      res_0_sum <= res_0_sum + score_0_x306;
      res_1_sum <= res_1_sum + score_1_x306;
      res_2_sum <= res_2_sum + score_2_x306;
      res_3_sum <= res_3_sum + score_3_x306;
      res_4_sum <= res_4_sum + score_4_x306;
      res_5_sum <= res_5_sum + score_5_x306;
      res_6_sum <= res_6_sum + score_6_x306;
      res_7_sum <= res_7_sum + score_7_x306;
      res_8_sum <= res_8_sum + score_8_x306;
      res_9_sum <= res_9_sum + score_9_x306;
   end
   else if(res_done_x307) begin
      res_0_sum <= res_0_sum + score_0_x307;
      res_1_sum <= res_1_sum + score_1_x307;
      res_2_sum <= res_2_sum + score_2_x307;
      res_3_sum <= res_3_sum + score_3_x307;
      res_4_sum <= res_4_sum + score_4_x307;
      res_5_sum <= res_5_sum + score_5_x307;
      res_6_sum <= res_6_sum + score_6_x307;
      res_7_sum <= res_7_sum + score_7_x307;
      res_8_sum <= res_8_sum + score_8_x307;
      res_9_sum <= res_9_sum + score_9_x307;
   end
   else if(res_done_x308) begin
      res_0_sum <= res_0_sum + score_0_x308;
      res_1_sum <= res_1_sum + score_1_x308;
      res_2_sum <= res_2_sum + score_2_x308;
      res_3_sum <= res_3_sum + score_3_x308;
      res_4_sum <= res_4_sum + score_4_x308;
      res_5_sum <= res_5_sum + score_5_x308;
      res_6_sum <= res_6_sum + score_6_x308;
      res_7_sum <= res_7_sum + score_7_x308;
      res_8_sum <= res_8_sum + score_8_x308;
      res_9_sum <= res_9_sum + score_9_x308;
   end
   else if(res_done_x309) begin
      res_0_sum <= res_0_sum + score_0_x309;
      res_1_sum <= res_1_sum + score_1_x309;
      res_2_sum <= res_2_sum + score_2_x309;
      res_3_sum <= res_3_sum + score_3_x309;
      res_4_sum <= res_4_sum + score_4_x309;
      res_5_sum <= res_5_sum + score_5_x309;
      res_6_sum <= res_6_sum + score_6_x309;
      res_7_sum <= res_7_sum + score_7_x309;
      res_8_sum <= res_8_sum + score_8_x309;
      res_9_sum <= res_9_sum + score_9_x309;
   end
   else if(res_done_x310) begin
      res_0_sum <= res_0_sum + score_0_x310;
      res_1_sum <= res_1_sum + score_1_x310;
      res_2_sum <= res_2_sum + score_2_x310;
      res_3_sum <= res_3_sum + score_3_x310;
      res_4_sum <= res_4_sum + score_4_x310;
      res_5_sum <= res_5_sum + score_5_x310;
      res_6_sum <= res_6_sum + score_6_x310;
      res_7_sum <= res_7_sum + score_7_x310;
      res_8_sum <= res_8_sum + score_8_x310;
      res_9_sum <= res_9_sum + score_9_x310;
   end
   else if(res_done_x311) begin
      res_0_sum <= res_0_sum + score_0_x311;
      res_1_sum <= res_1_sum + score_1_x311;
      res_2_sum <= res_2_sum + score_2_x311;
      res_3_sum <= res_3_sum + score_3_x311;
      res_4_sum <= res_4_sum + score_4_x311;
      res_5_sum <= res_5_sum + score_5_x311;
      res_6_sum <= res_6_sum + score_6_x311;
      res_7_sum <= res_7_sum + score_7_x311;
      res_8_sum <= res_8_sum + score_8_x311;
      res_9_sum <= res_9_sum + score_9_x311;
   end
   else if(res_done_x312) begin
      res_0_sum <= res_0_sum + score_0_x312;
      res_1_sum <= res_1_sum + score_1_x312;
      res_2_sum <= res_2_sum + score_2_x312;
      res_3_sum <= res_3_sum + score_3_x312;
      res_4_sum <= res_4_sum + score_4_x312;
      res_5_sum <= res_5_sum + score_5_x312;
      res_6_sum <= res_6_sum + score_6_x312;
      res_7_sum <= res_7_sum + score_7_x312;
      res_8_sum <= res_8_sum + score_8_x312;
      res_9_sum <= res_9_sum + score_9_x312;
   end
   else if(res_done_x313) begin
      res_0_sum <= res_0_sum + score_0_x313;
      res_1_sum <= res_1_sum + score_1_x313;
      res_2_sum <= res_2_sum + score_2_x313;
      res_3_sum <= res_3_sum + score_3_x313;
      res_4_sum <= res_4_sum + score_4_x313;
      res_5_sum <= res_5_sum + score_5_x313;
      res_6_sum <= res_6_sum + score_6_x313;
      res_7_sum <= res_7_sum + score_7_x313;
      res_8_sum <= res_8_sum + score_8_x313;
      res_9_sum <= res_9_sum + score_9_x313;
   end
   else if(res_done_x314) begin
      res_0_sum <= res_0_sum + score_0_x314;
      res_1_sum <= res_1_sum + score_1_x314;
      res_2_sum <= res_2_sum + score_2_x314;
      res_3_sum <= res_3_sum + score_3_x314;
      res_4_sum <= res_4_sum + score_4_x314;
      res_5_sum <= res_5_sum + score_5_x314;
      res_6_sum <= res_6_sum + score_6_x314;
      res_7_sum <= res_7_sum + score_7_x314;
      res_8_sum <= res_8_sum + score_8_x314;
      res_9_sum <= res_9_sum + score_9_x314;
   end
   else if(res_done_x315) begin
      res_0_sum <= res_0_sum + score_0_x315;
      res_1_sum <= res_1_sum + score_1_x315;
      res_2_sum <= res_2_sum + score_2_x315;
      res_3_sum <= res_3_sum + score_3_x315;
      res_4_sum <= res_4_sum + score_4_x315;
      res_5_sum <= res_5_sum + score_5_x315;
      res_6_sum <= res_6_sum + score_6_x315;
      res_7_sum <= res_7_sum + score_7_x315;
      res_8_sum <= res_8_sum + score_8_x315;
      res_9_sum <= res_9_sum + score_9_x315;
   end
   else if(res_done_x316) begin
      res_0_sum <= res_0_sum + score_0_x316;
      res_1_sum <= res_1_sum + score_1_x316;
      res_2_sum <= res_2_sum + score_2_x316;
      res_3_sum <= res_3_sum + score_3_x316;
      res_4_sum <= res_4_sum + score_4_x316;
      res_5_sum <= res_5_sum + score_5_x316;
      res_6_sum <= res_6_sum + score_6_x316;
      res_7_sum <= res_7_sum + score_7_x316;
      res_8_sum <= res_8_sum + score_8_x316;
      res_9_sum <= res_9_sum + score_9_x316;
   end
   else if(res_done_x317) begin
      res_0_sum <= res_0_sum + score_0_x317;
      res_1_sum <= res_1_sum + score_1_x317;
      res_2_sum <= res_2_sum + score_2_x317;
      res_3_sum <= res_3_sum + score_3_x317;
      res_4_sum <= res_4_sum + score_4_x317;
      res_5_sum <= res_5_sum + score_5_x317;
      res_6_sum <= res_6_sum + score_6_x317;
      res_7_sum <= res_7_sum + score_7_x317;
      res_8_sum <= res_8_sum + score_8_x317;
      res_9_sum <= res_9_sum + score_9_x317;
   end
   else if(res_done_x318) begin
      res_0_sum <= res_0_sum + score_0_x318;
      res_1_sum <= res_1_sum + score_1_x318;
      res_2_sum <= res_2_sum + score_2_x318;
      res_3_sum <= res_3_sum + score_3_x318;
      res_4_sum <= res_4_sum + score_4_x318;
      res_5_sum <= res_5_sum + score_5_x318;
      res_6_sum <= res_6_sum + score_6_x318;
      res_7_sum <= res_7_sum + score_7_x318;
      res_8_sum <= res_8_sum + score_8_x318;
      res_9_sum <= res_9_sum + score_9_x318;
   end
   else if(res_done_x319) begin
      res_0_sum <= res_0_sum + score_0_x319;
      res_1_sum <= res_1_sum + score_1_x319;
      res_2_sum <= res_2_sum + score_2_x319;
      res_3_sum <= res_3_sum + score_3_x319;
      res_4_sum <= res_4_sum + score_4_x319;
      res_5_sum <= res_5_sum + score_5_x319;
      res_6_sum <= res_6_sum + score_6_x319;
      res_7_sum <= res_7_sum + score_7_x319;
      res_8_sum <= res_8_sum + score_8_x319;
      res_9_sum <= res_9_sum + score_9_x319;
   end
   else if(res_done_x320) begin
      res_0_sum <= res_0_sum + score_0_x320;
      res_1_sum <= res_1_sum + score_1_x320;
      res_2_sum <= res_2_sum + score_2_x320;
      res_3_sum <= res_3_sum + score_3_x320;
      res_4_sum <= res_4_sum + score_4_x320;
      res_5_sum <= res_5_sum + score_5_x320;
      res_6_sum <= res_6_sum + score_6_x320;
      res_7_sum <= res_7_sum + score_7_x320;
      res_8_sum <= res_8_sum + score_8_x320;
      res_9_sum <= res_9_sum + score_9_x320;
   end
   else if(res_done_x321) begin
      res_0_sum <= res_0_sum + score_0_x321;
      res_1_sum <= res_1_sum + score_1_x321;
      res_2_sum <= res_2_sum + score_2_x321;
      res_3_sum <= res_3_sum + score_3_x321;
      res_4_sum <= res_4_sum + score_4_x321;
      res_5_sum <= res_5_sum + score_5_x321;
      res_6_sum <= res_6_sum + score_6_x321;
      res_7_sum <= res_7_sum + score_7_x321;
      res_8_sum <= res_8_sum + score_8_x321;
      res_9_sum <= res_9_sum + score_9_x321;
   end
   else if(res_done_x322) begin
      res_0_sum <= res_0_sum + score_0_x322;
      res_1_sum <= res_1_sum + score_1_x322;
      res_2_sum <= res_2_sum + score_2_x322;
      res_3_sum <= res_3_sum + score_3_x322;
      res_4_sum <= res_4_sum + score_4_x322;
      res_5_sum <= res_5_sum + score_5_x322;
      res_6_sum <= res_6_sum + score_6_x322;
      res_7_sum <= res_7_sum + score_7_x322;
      res_8_sum <= res_8_sum + score_8_x322;
      res_9_sum <= res_9_sum + score_9_x322;
   end
   else if(res_done_x323) begin
      res_0_sum <= res_0_sum + score_0_x323;
      res_1_sum <= res_1_sum + score_1_x323;
      res_2_sum <= res_2_sum + score_2_x323;
      res_3_sum <= res_3_sum + score_3_x323;
      res_4_sum <= res_4_sum + score_4_x323;
      res_5_sum <= res_5_sum + score_5_x323;
      res_6_sum <= res_6_sum + score_6_x323;
      res_7_sum <= res_7_sum + score_7_x323;
      res_8_sum <= res_8_sum + score_8_x323;
      res_9_sum <= res_9_sum + score_9_x323;
   end
   else if(res_done_x324) begin
      res_0_sum <= res_0_sum + score_0_x324;
      res_1_sum <= res_1_sum + score_1_x324;
      res_2_sum <= res_2_sum + score_2_x324;
      res_3_sum <= res_3_sum + score_3_x324;
      res_4_sum <= res_4_sum + score_4_x324;
      res_5_sum <= res_5_sum + score_5_x324;
      res_6_sum <= res_6_sum + score_6_x324;
      res_7_sum <= res_7_sum + score_7_x324;
      res_8_sum <= res_8_sum + score_8_x324;
      res_9_sum <= res_9_sum + score_9_x324;
   end
   else if(res_done_x325) begin
      res_0_sum <= res_0_sum + score_0_x325;
      res_1_sum <= res_1_sum + score_1_x325;
      res_2_sum <= res_2_sum + score_2_x325;
      res_3_sum <= res_3_sum + score_3_x325;
      res_4_sum <= res_4_sum + score_4_x325;
      res_5_sum <= res_5_sum + score_5_x325;
      res_6_sum <= res_6_sum + score_6_x325;
      res_7_sum <= res_7_sum + score_7_x325;
      res_8_sum <= res_8_sum + score_8_x325;
      res_9_sum <= res_9_sum + score_9_x325;
   end
   else if(res_done_x326) begin
      res_0_sum <= res_0_sum + score_0_x326;
      res_1_sum <= res_1_sum + score_1_x326;
      res_2_sum <= res_2_sum + score_2_x326;
      res_3_sum <= res_3_sum + score_3_x326;
      res_4_sum <= res_4_sum + score_4_x326;
      res_5_sum <= res_5_sum + score_5_x326;
      res_6_sum <= res_6_sum + score_6_x326;
      res_7_sum <= res_7_sum + score_7_x326;
      res_8_sum <= res_8_sum + score_8_x326;
      res_9_sum <= res_9_sum + score_9_x326;
   end
   else if(res_done_x327) begin
      res_0_sum <= res_0_sum + score_0_x327;
      res_1_sum <= res_1_sum + score_1_x327;
      res_2_sum <= res_2_sum + score_2_x327;
      res_3_sum <= res_3_sum + score_3_x327;
      res_4_sum <= res_4_sum + score_4_x327;
      res_5_sum <= res_5_sum + score_5_x327;
      res_6_sum <= res_6_sum + score_6_x327;
      res_7_sum <= res_7_sum + score_7_x327;
      res_8_sum <= res_8_sum + score_8_x327;
      res_9_sum <= res_9_sum + score_9_x327;
   end
   else if(res_done_x328) begin
      res_0_sum <= res_0_sum + score_0_x328;
      res_1_sum <= res_1_sum + score_1_x328;
      res_2_sum <= res_2_sum + score_2_x328;
      res_3_sum <= res_3_sum + score_3_x328;
      res_4_sum <= res_4_sum + score_4_x328;
      res_5_sum <= res_5_sum + score_5_x328;
      res_6_sum <= res_6_sum + score_6_x328;
      res_7_sum <= res_7_sum + score_7_x328;
      res_8_sum <= res_8_sum + score_8_x328;
      res_9_sum <= res_9_sum + score_9_x328;
   end
   else if(res_done_x329) begin
      res_0_sum <= res_0_sum + score_0_x329;
      res_1_sum <= res_1_sum + score_1_x329;
      res_2_sum <= res_2_sum + score_2_x329;
      res_3_sum <= res_3_sum + score_3_x329;
      res_4_sum <= res_4_sum + score_4_x329;
      res_5_sum <= res_5_sum + score_5_x329;
      res_6_sum <= res_6_sum + score_6_x329;
      res_7_sum <= res_7_sum + score_7_x329;
      res_8_sum <= res_8_sum + score_8_x329;
      res_9_sum <= res_9_sum + score_9_x329;
   end
   else if(res_done_x330) begin
      res_0_sum <= res_0_sum + score_0_x330;
      res_1_sum <= res_1_sum + score_1_x330;
      res_2_sum <= res_2_sum + score_2_x330;
      res_3_sum <= res_3_sum + score_3_x330;
      res_4_sum <= res_4_sum + score_4_x330;
      res_5_sum <= res_5_sum + score_5_x330;
      res_6_sum <= res_6_sum + score_6_x330;
      res_7_sum <= res_7_sum + score_7_x330;
      res_8_sum <= res_8_sum + score_8_x330;
      res_9_sum <= res_9_sum + score_9_x330;
   end
   else if(res_done_x331) begin
      res_0_sum <= res_0_sum + score_0_x331;
      res_1_sum <= res_1_sum + score_1_x331;
      res_2_sum <= res_2_sum + score_2_x331;
      res_3_sum <= res_3_sum + score_3_x331;
      res_4_sum <= res_4_sum + score_4_x331;
      res_5_sum <= res_5_sum + score_5_x331;
      res_6_sum <= res_6_sum + score_6_x331;
      res_7_sum <= res_7_sum + score_7_x331;
      res_8_sum <= res_8_sum + score_8_x331;
      res_9_sum <= res_9_sum + score_9_x331;
   end
   else if(res_done_x332) begin
      res_0_sum <= res_0_sum + score_0_x332;
      res_1_sum <= res_1_sum + score_1_x332;
      res_2_sum <= res_2_sum + score_2_x332;
      res_3_sum <= res_3_sum + score_3_x332;
      res_4_sum <= res_4_sum + score_4_x332;
      res_5_sum <= res_5_sum + score_5_x332;
      res_6_sum <= res_6_sum + score_6_x332;
      res_7_sum <= res_7_sum + score_7_x332;
      res_8_sum <= res_8_sum + score_8_x332;
      res_9_sum <= res_9_sum + score_9_x332;
   end
   else if(res_done_x333) begin
      res_0_sum <= res_0_sum + score_0_x333;
      res_1_sum <= res_1_sum + score_1_x333;
      res_2_sum <= res_2_sum + score_2_x333;
      res_3_sum <= res_3_sum + score_3_x333;
      res_4_sum <= res_4_sum + score_4_x333;
      res_5_sum <= res_5_sum + score_5_x333;
      res_6_sum <= res_6_sum + score_6_x333;
      res_7_sum <= res_7_sum + score_7_x333;
      res_8_sum <= res_8_sum + score_8_x333;
      res_9_sum <= res_9_sum + score_9_x333;
   end
   else if(res_done_x334) begin
      res_0_sum <= res_0_sum + score_0_x334;
      res_1_sum <= res_1_sum + score_1_x334;
      res_2_sum <= res_2_sum + score_2_x334;
      res_3_sum <= res_3_sum + score_3_x334;
      res_4_sum <= res_4_sum + score_4_x334;
      res_5_sum <= res_5_sum + score_5_x334;
      res_6_sum <= res_6_sum + score_6_x334;
      res_7_sum <= res_7_sum + score_7_x334;
      res_8_sum <= res_8_sum + score_8_x334;
      res_9_sum <= res_9_sum + score_9_x334;
   end
   else if(res_done_x335) begin
      res_0_sum <= res_0_sum + score_0_x335;
      res_1_sum <= res_1_sum + score_1_x335;
      res_2_sum <= res_2_sum + score_2_x335;
      res_3_sum <= res_3_sum + score_3_x335;
      res_4_sum <= res_4_sum + score_4_x335;
      res_5_sum <= res_5_sum + score_5_x335;
      res_6_sum <= res_6_sum + score_6_x335;
      res_7_sum <= res_7_sum + score_7_x335;
      res_8_sum <= res_8_sum + score_8_x335;
      res_9_sum <= res_9_sum + score_9_x335;
   end
   else if(res_done_x336) begin
      res_0_sum <= res_0_sum + score_0_x336;
      res_1_sum <= res_1_sum + score_1_x336;
      res_2_sum <= res_2_sum + score_2_x336;
      res_3_sum <= res_3_sum + score_3_x336;
      res_4_sum <= res_4_sum + score_4_x336;
      res_5_sum <= res_5_sum + score_5_x336;
      res_6_sum <= res_6_sum + score_6_x336;
      res_7_sum <= res_7_sum + score_7_x336;
      res_8_sum <= res_8_sum + score_8_x336;
      res_9_sum <= res_9_sum + score_9_x336;
   end
   else if(res_done_x337) begin
      res_0_sum <= res_0_sum + score_0_x337;
      res_1_sum <= res_1_sum + score_1_x337;
      res_2_sum <= res_2_sum + score_2_x337;
      res_3_sum <= res_3_sum + score_3_x337;
      res_4_sum <= res_4_sum + score_4_x337;
      res_5_sum <= res_5_sum + score_5_x337;
      res_6_sum <= res_6_sum + score_6_x337;
      res_7_sum <= res_7_sum + score_7_x337;
      res_8_sum <= res_8_sum + score_8_x337;
      res_9_sum <= res_9_sum + score_9_x337;
   end
   else if(res_done_x338) begin
      res_0_sum <= res_0_sum + score_0_x338;
      res_1_sum <= res_1_sum + score_1_x338;
      res_2_sum <= res_2_sum + score_2_x338;
      res_3_sum <= res_3_sum + score_3_x338;
      res_4_sum <= res_4_sum + score_4_x338;
      res_5_sum <= res_5_sum + score_5_x338;
      res_6_sum <= res_6_sum + score_6_x338;
      res_7_sum <= res_7_sum + score_7_x338;
      res_8_sum <= res_8_sum + score_8_x338;
      res_9_sum <= res_9_sum + score_9_x338;
   end
   else if(res_done_x339) begin
      res_0_sum <= res_0_sum + score_0_x339;
      res_1_sum <= res_1_sum + score_1_x339;
      res_2_sum <= res_2_sum + score_2_x339;
      res_3_sum <= res_3_sum + score_3_x339;
      res_4_sum <= res_4_sum + score_4_x339;
      res_5_sum <= res_5_sum + score_5_x339;
      res_6_sum <= res_6_sum + score_6_x339;
      res_7_sum <= res_7_sum + score_7_x339;
      res_8_sum <= res_8_sum + score_8_x339;
      res_9_sum <= res_9_sum + score_9_x339;
   end
   else if(res_done_x340) begin
      res_0_sum <= res_0_sum + score_0_x340;
      res_1_sum <= res_1_sum + score_1_x340;
      res_2_sum <= res_2_sum + score_2_x340;
      res_3_sum <= res_3_sum + score_3_x340;
      res_4_sum <= res_4_sum + score_4_x340;
      res_5_sum <= res_5_sum + score_5_x340;
      res_6_sum <= res_6_sum + score_6_x340;
      res_7_sum <= res_7_sum + score_7_x340;
      res_8_sum <= res_8_sum + score_8_x340;
      res_9_sum <= res_9_sum + score_9_x340;
   end
   else if(res_done_x341) begin
      res_0_sum <= res_0_sum + score_0_x341;
      res_1_sum <= res_1_sum + score_1_x341;
      res_2_sum <= res_2_sum + score_2_x341;
      res_3_sum <= res_3_sum + score_3_x341;
      res_4_sum <= res_4_sum + score_4_x341;
      res_5_sum <= res_5_sum + score_5_x341;
      res_6_sum <= res_6_sum + score_6_x341;
      res_7_sum <= res_7_sum + score_7_x341;
      res_8_sum <= res_8_sum + score_8_x341;
      res_9_sum <= res_9_sum + score_9_x341;
   end
   else if(res_done_x342) begin
      res_0_sum <= res_0_sum + score_0_x342;
      res_1_sum <= res_1_sum + score_1_x342;
      res_2_sum <= res_2_sum + score_2_x342;
      res_3_sum <= res_3_sum + score_3_x342;
      res_4_sum <= res_4_sum + score_4_x342;
      res_5_sum <= res_5_sum + score_5_x342;
      res_6_sum <= res_6_sum + score_6_x342;
      res_7_sum <= res_7_sum + score_7_x342;
      res_8_sum <= res_8_sum + score_8_x342;
      res_9_sum <= res_9_sum + score_9_x342;
   end
   else if(res_done_x343) begin
      res_0_sum <= res_0_sum + score_0_x343;
      res_1_sum <= res_1_sum + score_1_x343;
      res_2_sum <= res_2_sum + score_2_x343;
      res_3_sum <= res_3_sum + score_3_x343;
      res_4_sum <= res_4_sum + score_4_x343;
      res_5_sum <= res_5_sum + score_5_x343;
      res_6_sum <= res_6_sum + score_6_x343;
      res_7_sum <= res_7_sum + score_7_x343;
      res_8_sum <= res_8_sum + score_8_x343;
      res_9_sum <= res_9_sum + score_9_x343;
   end
   else if(res_done_x344) begin
      res_0_sum <= res_0_sum + score_0_x344;
      res_1_sum <= res_1_sum + score_1_x344;
      res_2_sum <= res_2_sum + score_2_x344;
      res_3_sum <= res_3_sum + score_3_x344;
      res_4_sum <= res_4_sum + score_4_x344;
      res_5_sum <= res_5_sum + score_5_x344;
      res_6_sum <= res_6_sum + score_6_x344;
      res_7_sum <= res_7_sum + score_7_x344;
      res_8_sum <= res_8_sum + score_8_x344;
      res_9_sum <= res_9_sum + score_9_x344;
   end
   else if(res_done_x345) begin
      res_0_sum <= res_0_sum + score_0_x345;
      res_1_sum <= res_1_sum + score_1_x345;
      res_2_sum <= res_2_sum + score_2_x345;
      res_3_sum <= res_3_sum + score_3_x345;
      res_4_sum <= res_4_sum + score_4_x345;
      res_5_sum <= res_5_sum + score_5_x345;
      res_6_sum <= res_6_sum + score_6_x345;
      res_7_sum <= res_7_sum + score_7_x345;
      res_8_sum <= res_8_sum + score_8_x345;
      res_9_sum <= res_9_sum + score_9_x345;
   end
   else if(res_done_x346) begin
      res_0_sum <= res_0_sum + score_0_x346;
      res_1_sum <= res_1_sum + score_1_x346;
      res_2_sum <= res_2_sum + score_2_x346;
      res_3_sum <= res_3_sum + score_3_x346;
      res_4_sum <= res_4_sum + score_4_x346;
      res_5_sum <= res_5_sum + score_5_x346;
      res_6_sum <= res_6_sum + score_6_x346;
      res_7_sum <= res_7_sum + score_7_x346;
      res_8_sum <= res_8_sum + score_8_x346;
      res_9_sum <= res_9_sum + score_9_x346;
   end
   else if(res_done_x347) begin
      res_0_sum <= res_0_sum + score_0_x347;
      res_1_sum <= res_1_sum + score_1_x347;
      res_2_sum <= res_2_sum + score_2_x347;
      res_3_sum <= res_3_sum + score_3_x347;
      res_4_sum <= res_4_sum + score_4_x347;
      res_5_sum <= res_5_sum + score_5_x347;
      res_6_sum <= res_6_sum + score_6_x347;
      res_7_sum <= res_7_sum + score_7_x347;
      res_8_sum <= res_8_sum + score_8_x347;
      res_9_sum <= res_9_sum + score_9_x347;
   end
   else if(res_done_x348) begin
      res_0_sum <= res_0_sum + score_0_x348;
      res_1_sum <= res_1_sum + score_1_x348;
      res_2_sum <= res_2_sum + score_2_x348;
      res_3_sum <= res_3_sum + score_3_x348;
      res_4_sum <= res_4_sum + score_4_x348;
      res_5_sum <= res_5_sum + score_5_x348;
      res_6_sum <= res_6_sum + score_6_x348;
      res_7_sum <= res_7_sum + score_7_x348;
      res_8_sum <= res_8_sum + score_8_x348;
      res_9_sum <= res_9_sum + score_9_x348;
   end
   else if(res_done_x349) begin
      res_0_sum <= res_0_sum + score_0_x349;
      res_1_sum <= res_1_sum + score_1_x349;
      res_2_sum <= res_2_sum + score_2_x349;
      res_3_sum <= res_3_sum + score_3_x349;
      res_4_sum <= res_4_sum + score_4_x349;
      res_5_sum <= res_5_sum + score_5_x349;
      res_6_sum <= res_6_sum + score_6_x349;
      res_7_sum <= res_7_sum + score_7_x349;
      res_8_sum <= res_8_sum + score_8_x349;
      res_9_sum <= res_9_sum + score_9_x349;
   end
   else if(res_done_x350) begin
      res_0_sum <= res_0_sum + score_0_x350;
      res_1_sum <= res_1_sum + score_1_x350;
      res_2_sum <= res_2_sum + score_2_x350;
      res_3_sum <= res_3_sum + score_3_x350;
      res_4_sum <= res_4_sum + score_4_x350;
      res_5_sum <= res_5_sum + score_5_x350;
      res_6_sum <= res_6_sum + score_6_x350;
      res_7_sum <= res_7_sum + score_7_x350;
      res_8_sum <= res_8_sum + score_8_x350;
      res_9_sum <= res_9_sum + score_9_x350;
   end
   else if(res_done_x351) begin
      res_0_sum <= res_0_sum + score_0_x351;
      res_1_sum <= res_1_sum + score_1_x351;
      res_2_sum <= res_2_sum + score_2_x351;
      res_3_sum <= res_3_sum + score_3_x351;
      res_4_sum <= res_4_sum + score_4_x351;
      res_5_sum <= res_5_sum + score_5_x351;
      res_6_sum <= res_6_sum + score_6_x351;
      res_7_sum <= res_7_sum + score_7_x351;
      res_8_sum <= res_8_sum + score_8_x351;
      res_9_sum <= res_9_sum + score_9_x351;
   end
   else if(res_done_x352) begin
      res_0_sum <= res_0_sum + score_0_x352;
      res_1_sum <= res_1_sum + score_1_x352;
      res_2_sum <= res_2_sum + score_2_x352;
      res_3_sum <= res_3_sum + score_3_x352;
      res_4_sum <= res_4_sum + score_4_x352;
      res_5_sum <= res_5_sum + score_5_x352;
      res_6_sum <= res_6_sum + score_6_x352;
      res_7_sum <= res_7_sum + score_7_x352;
      res_8_sum <= res_8_sum + score_8_x352;
      res_9_sum <= res_9_sum + score_9_x352;
   end
   else if(res_done_x353) begin
      res_0_sum <= res_0_sum + score_0_x353;
      res_1_sum <= res_1_sum + score_1_x353;
      res_2_sum <= res_2_sum + score_2_x353;
      res_3_sum <= res_3_sum + score_3_x353;
      res_4_sum <= res_4_sum + score_4_x353;
      res_5_sum <= res_5_sum + score_5_x353;
      res_6_sum <= res_6_sum + score_6_x353;
      res_7_sum <= res_7_sum + score_7_x353;
      res_8_sum <= res_8_sum + score_8_x353;
      res_9_sum <= res_9_sum + score_9_x353;
   end
   else if(res_done_x354) begin
      res_0_sum <= res_0_sum + score_0_x354;
      res_1_sum <= res_1_sum + score_1_x354;
      res_2_sum <= res_2_sum + score_2_x354;
      res_3_sum <= res_3_sum + score_3_x354;
      res_4_sum <= res_4_sum + score_4_x354;
      res_5_sum <= res_5_sum + score_5_x354;
      res_6_sum <= res_6_sum + score_6_x354;
      res_7_sum <= res_7_sum + score_7_x354;
      res_8_sum <= res_8_sum + score_8_x354;
      res_9_sum <= res_9_sum + score_9_x354;
   end
   else if(res_done_x355) begin
      res_0_sum <= res_0_sum + score_0_x355;
      res_1_sum <= res_1_sum + score_1_x355;
      res_2_sum <= res_2_sum + score_2_x355;
      res_3_sum <= res_3_sum + score_3_x355;
      res_4_sum <= res_4_sum + score_4_x355;
      res_5_sum <= res_5_sum + score_5_x355;
      res_6_sum <= res_6_sum + score_6_x355;
      res_7_sum <= res_7_sum + score_7_x355;
      res_8_sum <= res_8_sum + score_8_x355;
      res_9_sum <= res_9_sum + score_9_x355;
   end
   else if(res_done_x356) begin
      res_0_sum <= res_0_sum + score_0_x356;
      res_1_sum <= res_1_sum + score_1_x356;
      res_2_sum <= res_2_sum + score_2_x356;
      res_3_sum <= res_3_sum + score_3_x356;
      res_4_sum <= res_4_sum + score_4_x356;
      res_5_sum <= res_5_sum + score_5_x356;
      res_6_sum <= res_6_sum + score_6_x356;
      res_7_sum <= res_7_sum + score_7_x356;
      res_8_sum <= res_8_sum + score_8_x356;
      res_9_sum <= res_9_sum + score_9_x356;
   end
   else if(res_done_x357) begin
      res_0_sum <= res_0_sum + score_0_x357;
      res_1_sum <= res_1_sum + score_1_x357;
      res_2_sum <= res_2_sum + score_2_x357;
      res_3_sum <= res_3_sum + score_3_x357;
      res_4_sum <= res_4_sum + score_4_x357;
      res_5_sum <= res_5_sum + score_5_x357;
      res_6_sum <= res_6_sum + score_6_x357;
      res_7_sum <= res_7_sum + score_7_x357;
      res_8_sum <= res_8_sum + score_8_x357;
      res_9_sum <= res_9_sum + score_9_x357;
   end
   else if(res_done_x358) begin
      res_0_sum <= res_0_sum + score_0_x358;
      res_1_sum <= res_1_sum + score_1_x358;
      res_2_sum <= res_2_sum + score_2_x358;
      res_3_sum <= res_3_sum + score_3_x358;
      res_4_sum <= res_4_sum + score_4_x358;
      res_5_sum <= res_5_sum + score_5_x358;
      res_6_sum <= res_6_sum + score_6_x358;
      res_7_sum <= res_7_sum + score_7_x358;
      res_8_sum <= res_8_sum + score_8_x358;
      res_9_sum <= res_9_sum + score_9_x358;
   end
   else if(res_done_x359) begin
      res_0_sum <= res_0_sum + score_0_x359;
      res_1_sum <= res_1_sum + score_1_x359;
      res_2_sum <= res_2_sum + score_2_x359;
      res_3_sum <= res_3_sum + score_3_x359;
      res_4_sum <= res_4_sum + score_4_x359;
      res_5_sum <= res_5_sum + score_5_x359;
      res_6_sum <= res_6_sum + score_6_x359;
      res_7_sum <= res_7_sum + score_7_x359;
      res_8_sum <= res_8_sum + score_8_x359;
      res_9_sum <= res_9_sum + score_9_x359;
   end
   else if(res_done_x360) begin
      res_0_sum <= res_0_sum + score_0_x360;
      res_1_sum <= res_1_sum + score_1_x360;
      res_2_sum <= res_2_sum + score_2_x360;
      res_3_sum <= res_3_sum + score_3_x360;
      res_4_sum <= res_4_sum + score_4_x360;
      res_5_sum <= res_5_sum + score_5_x360;
      res_6_sum <= res_6_sum + score_6_x360;
      res_7_sum <= res_7_sum + score_7_x360;
      res_8_sum <= res_8_sum + score_8_x360;
      res_9_sum <= res_9_sum + score_9_x360;
   end
   else if(res_done_x361) begin
      res_0_sum <= res_0_sum + score_0_x361;
      res_1_sum <= res_1_sum + score_1_x361;
      res_2_sum <= res_2_sum + score_2_x361;
      res_3_sum <= res_3_sum + score_3_x361;
      res_4_sum <= res_4_sum + score_4_x361;
      res_5_sum <= res_5_sum + score_5_x361;
      res_6_sum <= res_6_sum + score_6_x361;
      res_7_sum <= res_7_sum + score_7_x361;
      res_8_sum <= res_8_sum + score_8_x361;
      res_9_sum <= res_9_sum + score_9_x361;
   end
   else if(res_done_x362) begin
      res_0_sum <= res_0_sum + score_0_x362;
      res_1_sum <= res_1_sum + score_1_x362;
      res_2_sum <= res_2_sum + score_2_x362;
      res_3_sum <= res_3_sum + score_3_x362;
      res_4_sum <= res_4_sum + score_4_x362;
      res_5_sum <= res_5_sum + score_5_x362;
      res_6_sum <= res_6_sum + score_6_x362;
      res_7_sum <= res_7_sum + score_7_x362;
      res_8_sum <= res_8_sum + score_8_x362;
      res_9_sum <= res_9_sum + score_9_x362;
   end
   else if(res_done_x363) begin
      res_0_sum <= res_0_sum + score_0_x363;
      res_1_sum <= res_1_sum + score_1_x363;
      res_2_sum <= res_2_sum + score_2_x363;
      res_3_sum <= res_3_sum + score_3_x363;
      res_4_sum <= res_4_sum + score_4_x363;
      res_5_sum <= res_5_sum + score_5_x363;
      res_6_sum <= res_6_sum + score_6_x363;
      res_7_sum <= res_7_sum + score_7_x363;
      res_8_sum <= res_8_sum + score_8_x363;
      res_9_sum <= res_9_sum + score_9_x363;
   end
   else if(res_done_x364) begin
      res_0_sum <= res_0_sum + score_0_x364;
      res_1_sum <= res_1_sum + score_1_x364;
      res_2_sum <= res_2_sum + score_2_x364;
      res_3_sum <= res_3_sum + score_3_x364;
      res_4_sum <= res_4_sum + score_4_x364;
      res_5_sum <= res_5_sum + score_5_x364;
      res_6_sum <= res_6_sum + score_6_x364;
      res_7_sum <= res_7_sum + score_7_x364;
      res_8_sum <= res_8_sum + score_8_x364;
      res_9_sum <= res_9_sum + score_9_x364;
   end
   else if(res_done_x365) begin
      res_0_sum <= res_0_sum + score_0_x365;
      res_1_sum <= res_1_sum + score_1_x365;
      res_2_sum <= res_2_sum + score_2_x365;
      res_3_sum <= res_3_sum + score_3_x365;
      res_4_sum <= res_4_sum + score_4_x365;
      res_5_sum <= res_5_sum + score_5_x365;
      res_6_sum <= res_6_sum + score_6_x365;
      res_7_sum <= res_7_sum + score_7_x365;
      res_8_sum <= res_8_sum + score_8_x365;
      res_9_sum <= res_9_sum + score_9_x365;
   end
   else if(res_done_x366) begin
      res_0_sum <= res_0_sum + score_0_x366;
      res_1_sum <= res_1_sum + score_1_x366;
      res_2_sum <= res_2_sum + score_2_x366;
      res_3_sum <= res_3_sum + score_3_x366;
      res_4_sum <= res_4_sum + score_4_x366;
      res_5_sum <= res_5_sum + score_5_x366;
      res_6_sum <= res_6_sum + score_6_x366;
      res_7_sum <= res_7_sum + score_7_x366;
      res_8_sum <= res_8_sum + score_8_x366;
      res_9_sum <= res_9_sum + score_9_x366;
   end
   else if(res_done_x367) begin
      res_0_sum <= res_0_sum + score_0_x367;
      res_1_sum <= res_1_sum + score_1_x367;
      res_2_sum <= res_2_sum + score_2_x367;
      res_3_sum <= res_3_sum + score_3_x367;
      res_4_sum <= res_4_sum + score_4_x367;
      res_5_sum <= res_5_sum + score_5_x367;
      res_6_sum <= res_6_sum + score_6_x367;
      res_7_sum <= res_7_sum + score_7_x367;
      res_8_sum <= res_8_sum + score_8_x367;
      res_9_sum <= res_9_sum + score_9_x367;
   end
   else if(res_done_x368) begin
      res_0_sum <= res_0_sum + score_0_x368;
      res_1_sum <= res_1_sum + score_1_x368;
      res_2_sum <= res_2_sum + score_2_x368;
      res_3_sum <= res_3_sum + score_3_x368;
      res_4_sum <= res_4_sum + score_4_x368;
      res_5_sum <= res_5_sum + score_5_x368;
      res_6_sum <= res_6_sum + score_6_x368;
      res_7_sum <= res_7_sum + score_7_x368;
      res_8_sum <= res_8_sum + score_8_x368;
      res_9_sum <= res_9_sum + score_9_x368;
   end
   else if(res_done_x369) begin
      res_0_sum <= res_0_sum + score_0_x369;
      res_1_sum <= res_1_sum + score_1_x369;
      res_2_sum <= res_2_sum + score_2_x369;
      res_3_sum <= res_3_sum + score_3_x369;
      res_4_sum <= res_4_sum + score_4_x369;
      res_5_sum <= res_5_sum + score_5_x369;
      res_6_sum <= res_6_sum + score_6_x369;
      res_7_sum <= res_7_sum + score_7_x369;
      res_8_sum <= res_8_sum + score_8_x369;
      res_9_sum <= res_9_sum + score_9_x369;
   end
   else if(res_done_x370) begin
      res_0_sum <= res_0_sum + score_0_x370;
      res_1_sum <= res_1_sum + score_1_x370;
      res_2_sum <= res_2_sum + score_2_x370;
      res_3_sum <= res_3_sum + score_3_x370;
      res_4_sum <= res_4_sum + score_4_x370;
      res_5_sum <= res_5_sum + score_5_x370;
      res_6_sum <= res_6_sum + score_6_x370;
      res_7_sum <= res_7_sum + score_7_x370;
      res_8_sum <= res_8_sum + score_8_x370;
      res_9_sum <= res_9_sum + score_9_x370;
   end
   else if(res_done_x371) begin
      res_0_sum <= res_0_sum + score_0_x371;
      res_1_sum <= res_1_sum + score_1_x371;
      res_2_sum <= res_2_sum + score_2_x371;
      res_3_sum <= res_3_sum + score_3_x371;
      res_4_sum <= res_4_sum + score_4_x371;
      res_5_sum <= res_5_sum + score_5_x371;
      res_6_sum <= res_6_sum + score_6_x371;
      res_7_sum <= res_7_sum + score_7_x371;
      res_8_sum <= res_8_sum + score_8_x371;
      res_9_sum <= res_9_sum + score_9_x371;
   end
   else if(res_done_x372) begin
      res_0_sum <= res_0_sum + score_0_x372;
      res_1_sum <= res_1_sum + score_1_x372;
      res_2_sum <= res_2_sum + score_2_x372;
      res_3_sum <= res_3_sum + score_3_x372;
      res_4_sum <= res_4_sum + score_4_x372;
      res_5_sum <= res_5_sum + score_5_x372;
      res_6_sum <= res_6_sum + score_6_x372;
      res_7_sum <= res_7_sum + score_7_x372;
      res_8_sum <= res_8_sum + score_8_x372;
      res_9_sum <= res_9_sum + score_9_x372;
   end
   else if(res_done_x373) begin
      res_0_sum <= res_0_sum + score_0_x373;
      res_1_sum <= res_1_sum + score_1_x373;
      res_2_sum <= res_2_sum + score_2_x373;
      res_3_sum <= res_3_sum + score_3_x373;
      res_4_sum <= res_4_sum + score_4_x373;
      res_5_sum <= res_5_sum + score_5_x373;
      res_6_sum <= res_6_sum + score_6_x373;
      res_7_sum <= res_7_sum + score_7_x373;
      res_8_sum <= res_8_sum + score_8_x373;
      res_9_sum <= res_9_sum + score_9_x373;
   end
   else if(res_done_x374) begin
      res_0_sum <= res_0_sum + score_0_x374;
      res_1_sum <= res_1_sum + score_1_x374;
      res_2_sum <= res_2_sum + score_2_x374;
      res_3_sum <= res_3_sum + score_3_x374;
      res_4_sum <= res_4_sum + score_4_x374;
      res_5_sum <= res_5_sum + score_5_x374;
      res_6_sum <= res_6_sum + score_6_x374;
      res_7_sum <= res_7_sum + score_7_x374;
      res_8_sum <= res_8_sum + score_8_x374;
      res_9_sum <= res_9_sum + score_9_x374;
   end
   else if(res_done_x375) begin
      res_0_sum <= res_0_sum + score_0_x375;
      res_1_sum <= res_1_sum + score_1_x375;
      res_2_sum <= res_2_sum + score_2_x375;
      res_3_sum <= res_3_sum + score_3_x375;
      res_4_sum <= res_4_sum + score_4_x375;
      res_5_sum <= res_5_sum + score_5_x375;
      res_6_sum <= res_6_sum + score_6_x375;
      res_7_sum <= res_7_sum + score_7_x375;
      res_8_sum <= res_8_sum + score_8_x375;
      res_9_sum <= res_9_sum + score_9_x375;
   end
   else if(res_done_x376) begin
      res_0_sum <= res_0_sum + score_0_x376;
      res_1_sum <= res_1_sum + score_1_x376;
      res_2_sum <= res_2_sum + score_2_x376;
      res_3_sum <= res_3_sum + score_3_x376;
      res_4_sum <= res_4_sum + score_4_x376;
      res_5_sum <= res_5_sum + score_5_x376;
      res_6_sum <= res_6_sum + score_6_x376;
      res_7_sum <= res_7_sum + score_7_x376;
      res_8_sum <= res_8_sum + score_8_x376;
      res_9_sum <= res_9_sum + score_9_x376;
   end
   else if(res_done_x377) begin
      res_0_sum <= res_0_sum + score_0_x377;
      res_1_sum <= res_1_sum + score_1_x377;
      res_2_sum <= res_2_sum + score_2_x377;
      res_3_sum <= res_3_sum + score_3_x377;
      res_4_sum <= res_4_sum + score_4_x377;
      res_5_sum <= res_5_sum + score_5_x377;
      res_6_sum <= res_6_sum + score_6_x377;
      res_7_sum <= res_7_sum + score_7_x377;
      res_8_sum <= res_8_sum + score_8_x377;
      res_9_sum <= res_9_sum + score_9_x377;
   end
   else if(res_done_x378) begin
      res_0_sum <= res_0_sum + score_0_x378;
      res_1_sum <= res_1_sum + score_1_x378;
      res_2_sum <= res_2_sum + score_2_x378;
      res_3_sum <= res_3_sum + score_3_x378;
      res_4_sum <= res_4_sum + score_4_x378;
      res_5_sum <= res_5_sum + score_5_x378;
      res_6_sum <= res_6_sum + score_6_x378;
      res_7_sum <= res_7_sum + score_7_x378;
      res_8_sum <= res_8_sum + score_8_x378;
      res_9_sum <= res_9_sum + score_9_x378;
   end
   else if(res_done_x379) begin
      res_0_sum <= res_0_sum + score_0_x379;
      res_1_sum <= res_1_sum + score_1_x379;
      res_2_sum <= res_2_sum + score_2_x379;
      res_3_sum <= res_3_sum + score_3_x379;
      res_4_sum <= res_4_sum + score_4_x379;
      res_5_sum <= res_5_sum + score_5_x379;
      res_6_sum <= res_6_sum + score_6_x379;
      res_7_sum <= res_7_sum + score_7_x379;
      res_8_sum <= res_8_sum + score_8_x379;
      res_9_sum <= res_9_sum + score_9_x379;
   end
   else if(res_done_x380) begin
      res_0_sum <= res_0_sum + score_0_x380;
      res_1_sum <= res_1_sum + score_1_x380;
      res_2_sum <= res_2_sum + score_2_x380;
      res_3_sum <= res_3_sum + score_3_x380;
      res_4_sum <= res_4_sum + score_4_x380;
      res_5_sum <= res_5_sum + score_5_x380;
      res_6_sum <= res_6_sum + score_6_x380;
      res_7_sum <= res_7_sum + score_7_x380;
      res_8_sum <= res_8_sum + score_8_x380;
      res_9_sum <= res_9_sum + score_9_x380;
   end
   else if(res_done_x381) begin
      res_0_sum <= res_0_sum + score_0_x381;
      res_1_sum <= res_1_sum + score_1_x381;
      res_2_sum <= res_2_sum + score_2_x381;
      res_3_sum <= res_3_sum + score_3_x381;
      res_4_sum <= res_4_sum + score_4_x381;
      res_5_sum <= res_5_sum + score_5_x381;
      res_6_sum <= res_6_sum + score_6_x381;
      res_7_sum <= res_7_sum + score_7_x381;
      res_8_sum <= res_8_sum + score_8_x381;
      res_9_sum <= res_9_sum + score_9_x381;
   end
   else if(res_done_x382) begin
      res_0_sum <= res_0_sum + score_0_x382;
      res_1_sum <= res_1_sum + score_1_x382;
      res_2_sum <= res_2_sum + score_2_x382;
      res_3_sum <= res_3_sum + score_3_x382;
      res_4_sum <= res_4_sum + score_4_x382;
      res_5_sum <= res_5_sum + score_5_x382;
      res_6_sum <= res_6_sum + score_6_x382;
      res_7_sum <= res_7_sum + score_7_x382;
      res_8_sum <= res_8_sum + score_8_x382;
      res_9_sum <= res_9_sum + score_9_x382;
   end
   else if(res_done_x383) begin
      res_0_sum <= res_0_sum + score_0_x383;
      res_1_sum <= res_1_sum + score_1_x383;
      res_2_sum <= res_2_sum + score_2_x383;
      res_3_sum <= res_3_sum + score_3_x383;
      res_4_sum <= res_4_sum + score_4_x383;
      res_5_sum <= res_5_sum + score_5_x383;
      res_6_sum <= res_6_sum + score_6_x383;
      res_7_sum <= res_7_sum + score_7_x383;
      res_8_sum <= res_8_sum + score_8_x383;
      res_9_sum <= res_9_sum + score_9_x383;
   end
   else if(res_done_x384) begin
      res_0_sum <= res_0_sum + score_0_x384;
      res_1_sum <= res_1_sum + score_1_x384;
      res_2_sum <= res_2_sum + score_2_x384;
      res_3_sum <= res_3_sum + score_3_x384;
      res_4_sum <= res_4_sum + score_4_x384;
      res_5_sum <= res_5_sum + score_5_x384;
      res_6_sum <= res_6_sum + score_6_x384;
      res_7_sum <= res_7_sum + score_7_x384;
      res_8_sum <= res_8_sum + score_8_x384;
      res_9_sum <= res_9_sum + score_9_x384;
   end
   else if(res_done_x385) begin
      res_0_sum <= res_0_sum + score_0_x385;
      res_1_sum <= res_1_sum + score_1_x385;
      res_2_sum <= res_2_sum + score_2_x385;
      res_3_sum <= res_3_sum + score_3_x385;
      res_4_sum <= res_4_sum + score_4_x385;
      res_5_sum <= res_5_sum + score_5_x385;
      res_6_sum <= res_6_sum + score_6_x385;
      res_7_sum <= res_7_sum + score_7_x385;
      res_8_sum <= res_8_sum + score_8_x385;
      res_9_sum <= res_9_sum + score_9_x385;
   end
   else if(res_done_x386) begin
      res_0_sum <= res_0_sum + score_0_x386;
      res_1_sum <= res_1_sum + score_1_x386;
      res_2_sum <= res_2_sum + score_2_x386;
      res_3_sum <= res_3_sum + score_3_x386;
      res_4_sum <= res_4_sum + score_4_x386;
      res_5_sum <= res_5_sum + score_5_x386;
      res_6_sum <= res_6_sum + score_6_x386;
      res_7_sum <= res_7_sum + score_7_x386;
      res_8_sum <= res_8_sum + score_8_x386;
      res_9_sum <= res_9_sum + score_9_x386;
   end
   else if(res_done_x387) begin
      res_0_sum <= res_0_sum + score_0_x387;
      res_1_sum <= res_1_sum + score_1_x387;
      res_2_sum <= res_2_sum + score_2_x387;
      res_3_sum <= res_3_sum + score_3_x387;
      res_4_sum <= res_4_sum + score_4_x387;
      res_5_sum <= res_5_sum + score_5_x387;
      res_6_sum <= res_6_sum + score_6_x387;
      res_7_sum <= res_7_sum + score_7_x387;
      res_8_sum <= res_8_sum + score_8_x387;
      res_9_sum <= res_9_sum + score_9_x387;
   end
   else if(res_done_x388) begin
      res_0_sum <= res_0_sum + score_0_x388;
      res_1_sum <= res_1_sum + score_1_x388;
      res_2_sum <= res_2_sum + score_2_x388;
      res_3_sum <= res_3_sum + score_3_x388;
      res_4_sum <= res_4_sum + score_4_x388;
      res_5_sum <= res_5_sum + score_5_x388;
      res_6_sum <= res_6_sum + score_6_x388;
      res_7_sum <= res_7_sum + score_7_x388;
      res_8_sum <= res_8_sum + score_8_x388;
      res_9_sum <= res_9_sum + score_9_x388;
   end
   else if(res_done_x389) begin
      res_0_sum <= res_0_sum + score_0_x389;
      res_1_sum <= res_1_sum + score_1_x389;
      res_2_sum <= res_2_sum + score_2_x389;
      res_3_sum <= res_3_sum + score_3_x389;
      res_4_sum <= res_4_sum + score_4_x389;
      res_5_sum <= res_5_sum + score_5_x389;
      res_6_sum <= res_6_sum + score_6_x389;
      res_7_sum <= res_7_sum + score_7_x389;
      res_8_sum <= res_8_sum + score_8_x389;
      res_9_sum <= res_9_sum + score_9_x389;
   end
   else if(res_done_x390) begin
      res_0_sum <= res_0_sum + score_0_x390;
      res_1_sum <= res_1_sum + score_1_x390;
      res_2_sum <= res_2_sum + score_2_x390;
      res_3_sum <= res_3_sum + score_3_x390;
      res_4_sum <= res_4_sum + score_4_x390;
      res_5_sum <= res_5_sum + score_5_x390;
      res_6_sum <= res_6_sum + score_6_x390;
      res_7_sum <= res_7_sum + score_7_x390;
      res_8_sum <= res_8_sum + score_8_x390;
      res_9_sum <= res_9_sum + score_9_x390;
   end
   else if(res_done_x391) begin
      res_0_sum <= res_0_sum + score_0_x391;
      res_1_sum <= res_1_sum + score_1_x391;
      res_2_sum <= res_2_sum + score_2_x391;
      res_3_sum <= res_3_sum + score_3_x391;
      res_4_sum <= res_4_sum + score_4_x391;
      res_5_sum <= res_5_sum + score_5_x391;
      res_6_sum <= res_6_sum + score_6_x391;
      res_7_sum <= res_7_sum + score_7_x391;
      res_8_sum <= res_8_sum + score_8_x391;
      res_9_sum <= res_9_sum + score_9_x391;
   end
   else if(res_done_x392) begin
      res_0_sum <= res_0_sum + score_0_x392;
      res_1_sum <= res_1_sum + score_1_x392;
      res_2_sum <= res_2_sum + score_2_x392;
      res_3_sum <= res_3_sum + score_3_x392;
      res_4_sum <= res_4_sum + score_4_x392;
      res_5_sum <= res_5_sum + score_5_x392;
      res_6_sum <= res_6_sum + score_6_x392;
      res_7_sum <= res_7_sum + score_7_x392;
      res_8_sum <= res_8_sum + score_8_x392;
      res_9_sum <= res_9_sum + score_9_x392;
   end
   else if(res_done_x393) begin
      res_0_sum <= res_0_sum + score_0_x393;
      res_1_sum <= res_1_sum + score_1_x393;
      res_2_sum <= res_2_sum + score_2_x393;
      res_3_sum <= res_3_sum + score_3_x393;
      res_4_sum <= res_4_sum + score_4_x393;
      res_5_sum <= res_5_sum + score_5_x393;
      res_6_sum <= res_6_sum + score_6_x393;
      res_7_sum <= res_7_sum + score_7_x393;
      res_8_sum <= res_8_sum + score_8_x393;
      res_9_sum <= res_9_sum + score_9_x393;
   end
   else if(res_done_x394) begin
      res_0_sum <= res_0_sum + score_0_x394;
      res_1_sum <= res_1_sum + score_1_x394;
      res_2_sum <= res_2_sum + score_2_x394;
      res_3_sum <= res_3_sum + score_3_x394;
      res_4_sum <= res_4_sum + score_4_x394;
      res_5_sum <= res_5_sum + score_5_x394;
      res_6_sum <= res_6_sum + score_6_x394;
      res_7_sum <= res_7_sum + score_7_x394;
      res_8_sum <= res_8_sum + score_8_x394;
      res_9_sum <= res_9_sum + score_9_x394;
   end
   else if(res_done_x395) begin
      res_0_sum <= res_0_sum + score_0_x395;
      res_1_sum <= res_1_sum + score_1_x395;
      res_2_sum <= res_2_sum + score_2_x395;
      res_3_sum <= res_3_sum + score_3_x395;
      res_4_sum <= res_4_sum + score_4_x395;
      res_5_sum <= res_5_sum + score_5_x395;
      res_6_sum <= res_6_sum + score_6_x395;
      res_7_sum <= res_7_sum + score_7_x395;
      res_8_sum <= res_8_sum + score_8_x395;
      res_9_sum <= res_9_sum + score_9_x395;
   end
   else if(res_done_x396) begin
      res_0_sum <= res_0_sum + score_0_x396;
      res_1_sum <= res_1_sum + score_1_x396;
      res_2_sum <= res_2_sum + score_2_x396;
      res_3_sum <= res_3_sum + score_3_x396;
      res_4_sum <= res_4_sum + score_4_x396;
      res_5_sum <= res_5_sum + score_5_x396;
      res_6_sum <= res_6_sum + score_6_x396;
      res_7_sum <= res_7_sum + score_7_x396;
      res_8_sum <= res_8_sum + score_8_x396;
      res_9_sum <= res_9_sum + score_9_x396;
   end
   else if(res_done_x397) begin
      res_0_sum <= res_0_sum + score_0_x397;
      res_1_sum <= res_1_sum + score_1_x397;
      res_2_sum <= res_2_sum + score_2_x397;
      res_3_sum <= res_3_sum + score_3_x397;
      res_4_sum <= res_4_sum + score_4_x397;
      res_5_sum <= res_5_sum + score_5_x397;
      res_6_sum <= res_6_sum + score_6_x397;
      res_7_sum <= res_7_sum + score_7_x397;
      res_8_sum <= res_8_sum + score_8_x397;
      res_9_sum <= res_9_sum + score_9_x397;
   end
   else if(res_done_x398) begin
      res_0_sum <= res_0_sum + score_0_x398;
      res_1_sum <= res_1_sum + score_1_x398;
      res_2_sum <= res_2_sum + score_2_x398;
      res_3_sum <= res_3_sum + score_3_x398;
      res_4_sum <= res_4_sum + score_4_x398;
      res_5_sum <= res_5_sum + score_5_x398;
      res_6_sum <= res_6_sum + score_6_x398;
      res_7_sum <= res_7_sum + score_7_x398;
      res_8_sum <= res_8_sum + score_8_x398;
      res_9_sum <= res_9_sum + score_9_x398;
   end
   else if(res_done_x399) begin
      res_0_sum <= res_0_sum + score_0_x399;
      res_1_sum <= res_1_sum + score_1_x399;
      res_2_sum <= res_2_sum + score_2_x399;
      res_3_sum <= res_3_sum + score_3_x399;
      res_4_sum <= res_4_sum + score_4_x399;
      res_5_sum <= res_5_sum + score_5_x399;
      res_6_sum <= res_6_sum + score_6_x399;
      res_7_sum <= res_7_sum + score_7_x399;
      res_8_sum <= res_8_sum + score_8_x399;
      res_9_sum <= res_9_sum + score_9_x399;
   end
   else if(res_done_x400) begin
      res_0_sum <= res_0_sum + score_0_x400;
      res_1_sum <= res_1_sum + score_1_x400;
      res_2_sum <= res_2_sum + score_2_x400;
      res_3_sum <= res_3_sum + score_3_x400;
      res_4_sum <= res_4_sum + score_4_x400;
      res_5_sum <= res_5_sum + score_5_x400;
      res_6_sum <= res_6_sum + score_6_x400;
      res_7_sum <= res_7_sum + score_7_x400;
      res_8_sum <= res_8_sum + score_8_x400;
      res_9_sum <= res_9_sum + score_9_x400;
   end
   else if(res_done_x401) begin
      res_0_sum <= res_0_sum + score_0_x401;
      res_1_sum <= res_1_sum + score_1_x401;
      res_2_sum <= res_2_sum + score_2_x401;
      res_3_sum <= res_3_sum + score_3_x401;
      res_4_sum <= res_4_sum + score_4_x401;
      res_5_sum <= res_5_sum + score_5_x401;
      res_6_sum <= res_6_sum + score_6_x401;
      res_7_sum <= res_7_sum + score_7_x401;
      res_8_sum <= res_8_sum + score_8_x401;
      res_9_sum <= res_9_sum + score_9_x401;
   end
   else if(res_done_x402) begin
      res_0_sum <= res_0_sum + score_0_x402;
      res_1_sum <= res_1_sum + score_1_x402;
      res_2_sum <= res_2_sum + score_2_x402;
      res_3_sum <= res_3_sum + score_3_x402;
      res_4_sum <= res_4_sum + score_4_x402;
      res_5_sum <= res_5_sum + score_5_x402;
      res_6_sum <= res_6_sum + score_6_x402;
      res_7_sum <= res_7_sum + score_7_x402;
      res_8_sum <= res_8_sum + score_8_x402;
      res_9_sum <= res_9_sum + score_9_x402;
   end
   else if(res_done_x403) begin
      res_0_sum <= res_0_sum + score_0_x403;
      res_1_sum <= res_1_sum + score_1_x403;
      res_2_sum <= res_2_sum + score_2_x403;
      res_3_sum <= res_3_sum + score_3_x403;
      res_4_sum <= res_4_sum + score_4_x403;
      res_5_sum <= res_5_sum + score_5_x403;
      res_6_sum <= res_6_sum + score_6_x403;
      res_7_sum <= res_7_sum + score_7_x403;
      res_8_sum <= res_8_sum + score_8_x403;
      res_9_sum <= res_9_sum + score_9_x403;
   end
   else if(res_done_x404) begin
      res_0_sum <= res_0_sum + score_0_x404;
      res_1_sum <= res_1_sum + score_1_x404;
      res_2_sum <= res_2_sum + score_2_x404;
      res_3_sum <= res_3_sum + score_3_x404;
      res_4_sum <= res_4_sum + score_4_x404;
      res_5_sum <= res_5_sum + score_5_x404;
      res_6_sum <= res_6_sum + score_6_x404;
      res_7_sum <= res_7_sum + score_7_x404;
      res_8_sum <= res_8_sum + score_8_x404;
      res_9_sum <= res_9_sum + score_9_x404;
   end
   else if(res_done_x405) begin
      res_0_sum <= res_0_sum + score_0_x405;
      res_1_sum <= res_1_sum + score_1_x405;
      res_2_sum <= res_2_sum + score_2_x405;
      res_3_sum <= res_3_sum + score_3_x405;
      res_4_sum <= res_4_sum + score_4_x405;
      res_5_sum <= res_5_sum + score_5_x405;
      res_6_sum <= res_6_sum + score_6_x405;
      res_7_sum <= res_7_sum + score_7_x405;
      res_8_sum <= res_8_sum + score_8_x405;
      res_9_sum <= res_9_sum + score_9_x405;
   end
   else if(res_done_x406) begin
      res_0_sum <= res_0_sum + score_0_x406;
      res_1_sum <= res_1_sum + score_1_x406;
      res_2_sum <= res_2_sum + score_2_x406;
      res_3_sum <= res_3_sum + score_3_x406;
      res_4_sum <= res_4_sum + score_4_x406;
      res_5_sum <= res_5_sum + score_5_x406;
      res_6_sum <= res_6_sum + score_6_x406;
      res_7_sum <= res_7_sum + score_7_x406;
      res_8_sum <= res_8_sum + score_8_x406;
      res_9_sum <= res_9_sum + score_9_x406;
   end
   else if(res_done_x407) begin
      res_0_sum <= res_0_sum + score_0_x407;
      res_1_sum <= res_1_sum + score_1_x407;
      res_2_sum <= res_2_sum + score_2_x407;
      res_3_sum <= res_3_sum + score_3_x407;
      res_4_sum <= res_4_sum + score_4_x407;
      res_5_sum <= res_5_sum + score_5_x407;
      res_6_sum <= res_6_sum + score_6_x407;
      res_7_sum <= res_7_sum + score_7_x407;
      res_8_sum <= res_8_sum + score_8_x407;
      res_9_sum <= res_9_sum + score_9_x407;
   end
   else if(res_done_x408) begin
      res_0_sum <= res_0_sum + score_0_x408;
      res_1_sum <= res_1_sum + score_1_x408;
      res_2_sum <= res_2_sum + score_2_x408;
      res_3_sum <= res_3_sum + score_3_x408;
      res_4_sum <= res_4_sum + score_4_x408;
      res_5_sum <= res_5_sum + score_5_x408;
      res_6_sum <= res_6_sum + score_6_x408;
      res_7_sum <= res_7_sum + score_7_x408;
      res_8_sum <= res_8_sum + score_8_x408;
      res_9_sum <= res_9_sum + score_9_x408;
   end
   else if(res_done_x409) begin
      res_0_sum <= res_0_sum + score_0_x409;
      res_1_sum <= res_1_sum + score_1_x409;
      res_2_sum <= res_2_sum + score_2_x409;
      res_3_sum <= res_3_sum + score_3_x409;
      res_4_sum <= res_4_sum + score_4_x409;
      res_5_sum <= res_5_sum + score_5_x409;
      res_6_sum <= res_6_sum + score_6_x409;
      res_7_sum <= res_7_sum + score_7_x409;
      res_8_sum <= res_8_sum + score_8_x409;
      res_9_sum <= res_9_sum + score_9_x409;
   end
   else if(res_done_x410) begin
      res_0_sum <= res_0_sum + score_0_x410;
      res_1_sum <= res_1_sum + score_1_x410;
      res_2_sum <= res_2_sum + score_2_x410;
      res_3_sum <= res_3_sum + score_3_x410;
      res_4_sum <= res_4_sum + score_4_x410;
      res_5_sum <= res_5_sum + score_5_x410;
      res_6_sum <= res_6_sum + score_6_x410;
      res_7_sum <= res_7_sum + score_7_x410;
      res_8_sum <= res_8_sum + score_8_x410;
      res_9_sum <= res_9_sum + score_9_x410;
   end
   else if(res_done_x411) begin
      res_0_sum <= res_0_sum + score_0_x411;
      res_1_sum <= res_1_sum + score_1_x411;
      res_2_sum <= res_2_sum + score_2_x411;
      res_3_sum <= res_3_sum + score_3_x411;
      res_4_sum <= res_4_sum + score_4_x411;
      res_5_sum <= res_5_sum + score_5_x411;
      res_6_sum <= res_6_sum + score_6_x411;
      res_7_sum <= res_7_sum + score_7_x411;
      res_8_sum <= res_8_sum + score_8_x411;
      res_9_sum <= res_9_sum + score_9_x411;
   end
   else if(res_done_x412) begin
      res_0_sum <= res_0_sum + score_0_x412;
      res_1_sum <= res_1_sum + score_1_x412;
      res_2_sum <= res_2_sum + score_2_x412;
      res_3_sum <= res_3_sum + score_3_x412;
      res_4_sum <= res_4_sum + score_4_x412;
      res_5_sum <= res_5_sum + score_5_x412;
      res_6_sum <= res_6_sum + score_6_x412;
      res_7_sum <= res_7_sum + score_7_x412;
      res_8_sum <= res_8_sum + score_8_x412;
      res_9_sum <= res_9_sum + score_9_x412;
   end
   else if(res_done_x413) begin
      res_0_sum <= res_0_sum + score_0_x413;
      res_1_sum <= res_1_sum + score_1_x413;
      res_2_sum <= res_2_sum + score_2_x413;
      res_3_sum <= res_3_sum + score_3_x413;
      res_4_sum <= res_4_sum + score_4_x413;
      res_5_sum <= res_5_sum + score_5_x413;
      res_6_sum <= res_6_sum + score_6_x413;
      res_7_sum <= res_7_sum + score_7_x413;
      res_8_sum <= res_8_sum + score_8_x413;
      res_9_sum <= res_9_sum + score_9_x413;
   end
   else if(res_done_x414) begin
      res_0_sum <= res_0_sum + score_0_x414;
      res_1_sum <= res_1_sum + score_1_x414;
      res_2_sum <= res_2_sum + score_2_x414;
      res_3_sum <= res_3_sum + score_3_x414;
      res_4_sum <= res_4_sum + score_4_x414;
      res_5_sum <= res_5_sum + score_5_x414;
      res_6_sum <= res_6_sum + score_6_x414;
      res_7_sum <= res_7_sum + score_7_x414;
      res_8_sum <= res_8_sum + score_8_x414;
      res_9_sum <= res_9_sum + score_9_x414;
   end
   else if(res_done_x415) begin
      res_0_sum <= res_0_sum + score_0_x415;
      res_1_sum <= res_1_sum + score_1_x415;
      res_2_sum <= res_2_sum + score_2_x415;
      res_3_sum <= res_3_sum + score_3_x415;
      res_4_sum <= res_4_sum + score_4_x415;
      res_5_sum <= res_5_sum + score_5_x415;
      res_6_sum <= res_6_sum + score_6_x415;
      res_7_sum <= res_7_sum + score_7_x415;
      res_8_sum <= res_8_sum + score_8_x415;
      res_9_sum <= res_9_sum + score_9_x415;
   end
   else if(res_done_x416) begin
      res_0_sum <= res_0_sum + score_0_x416;
      res_1_sum <= res_1_sum + score_1_x416;
      res_2_sum <= res_2_sum + score_2_x416;
      res_3_sum <= res_3_sum + score_3_x416;
      res_4_sum <= res_4_sum + score_4_x416;
      res_5_sum <= res_5_sum + score_5_x416;
      res_6_sum <= res_6_sum + score_6_x416;
      res_7_sum <= res_7_sum + score_7_x416;
      res_8_sum <= res_8_sum + score_8_x416;
      res_9_sum <= res_9_sum + score_9_x416;
   end
   else if(res_done_x417) begin
      res_0_sum <= res_0_sum + score_0_x417;
      res_1_sum <= res_1_sum + score_1_x417;
      res_2_sum <= res_2_sum + score_2_x417;
      res_3_sum <= res_3_sum + score_3_x417;
      res_4_sum <= res_4_sum + score_4_x417;
      res_5_sum <= res_5_sum + score_5_x417;
      res_6_sum <= res_6_sum + score_6_x417;
      res_7_sum <= res_7_sum + score_7_x417;
      res_8_sum <= res_8_sum + score_8_x417;
      res_9_sum <= res_9_sum + score_9_x417;
   end
   else if(res_done_x418) begin
      res_0_sum <= res_0_sum + score_0_x418;
      res_1_sum <= res_1_sum + score_1_x418;
      res_2_sum <= res_2_sum + score_2_x418;
      res_3_sum <= res_3_sum + score_3_x418;
      res_4_sum <= res_4_sum + score_4_x418;
      res_5_sum <= res_5_sum + score_5_x418;
      res_6_sum <= res_6_sum + score_6_x418;
      res_7_sum <= res_7_sum + score_7_x418;
      res_8_sum <= res_8_sum + score_8_x418;
      res_9_sum <= res_9_sum + score_9_x418;
   end
   else if(res_done_x419) begin
      res_0_sum <= res_0_sum + score_0_x419;
      res_1_sum <= res_1_sum + score_1_x419;
      res_2_sum <= res_2_sum + score_2_x419;
      res_3_sum <= res_3_sum + score_3_x419;
      res_4_sum <= res_4_sum + score_4_x419;
      res_5_sum <= res_5_sum + score_5_x419;
      res_6_sum <= res_6_sum + score_6_x419;
      res_7_sum <= res_7_sum + score_7_x419;
      res_8_sum <= res_8_sum + score_8_x419;
      res_9_sum <= res_9_sum + score_9_x419;
   end
   else if(res_done_x420) begin
      res_0_sum <= res_0_sum + score_0_x420;
      res_1_sum <= res_1_sum + score_1_x420;
      res_2_sum <= res_2_sum + score_2_x420;
      res_3_sum <= res_3_sum + score_3_x420;
      res_4_sum <= res_4_sum + score_4_x420;
      res_5_sum <= res_5_sum + score_5_x420;
      res_6_sum <= res_6_sum + score_6_x420;
      res_7_sum <= res_7_sum + score_7_x420;
      res_8_sum <= res_8_sum + score_8_x420;
      res_9_sum <= res_9_sum + score_9_x420;
   end
   else if(res_done_x421) begin
      res_0_sum <= res_0_sum + score_0_x421;
      res_1_sum <= res_1_sum + score_1_x421;
      res_2_sum <= res_2_sum + score_2_x421;
      res_3_sum <= res_3_sum + score_3_x421;
      res_4_sum <= res_4_sum + score_4_x421;
      res_5_sum <= res_5_sum + score_5_x421;
      res_6_sum <= res_6_sum + score_6_x421;
      res_7_sum <= res_7_sum + score_7_x421;
      res_8_sum <= res_8_sum + score_8_x421;
      res_9_sum <= res_9_sum + score_9_x421;
   end
   else if(res_done_x422) begin
      res_0_sum <= res_0_sum + score_0_x422;
      res_1_sum <= res_1_sum + score_1_x422;
      res_2_sum <= res_2_sum + score_2_x422;
      res_3_sum <= res_3_sum + score_3_x422;
      res_4_sum <= res_4_sum + score_4_x422;
      res_5_sum <= res_5_sum + score_5_x422;
      res_6_sum <= res_6_sum + score_6_x422;
      res_7_sum <= res_7_sum + score_7_x422;
      res_8_sum <= res_8_sum + score_8_x422;
      res_9_sum <= res_9_sum + score_9_x422;
   end
   else if(res_done_x423) begin
      res_0_sum <= res_0_sum + score_0_x423;
      res_1_sum <= res_1_sum + score_1_x423;
      res_2_sum <= res_2_sum + score_2_x423;
      res_3_sum <= res_3_sum + score_3_x423;
      res_4_sum <= res_4_sum + score_4_x423;
      res_5_sum <= res_5_sum + score_5_x423;
      res_6_sum <= res_6_sum + score_6_x423;
      res_7_sum <= res_7_sum + score_7_x423;
      res_8_sum <= res_8_sum + score_8_x423;
      res_9_sum <= res_9_sum + score_9_x423;
   end
   else if(res_done_x424) begin
      res_0_sum <= res_0_sum + score_0_x424;
      res_1_sum <= res_1_sum + score_1_x424;
      res_2_sum <= res_2_sum + score_2_x424;
      res_3_sum <= res_3_sum + score_3_x424;
      res_4_sum <= res_4_sum + score_4_x424;
      res_5_sum <= res_5_sum + score_5_x424;
      res_6_sum <= res_6_sum + score_6_x424;
      res_7_sum <= res_7_sum + score_7_x424;
      res_8_sum <= res_8_sum + score_8_x424;
      res_9_sum <= res_9_sum + score_9_x424;
   end
   else if(res_done_x425) begin
      res_0_sum <= res_0_sum + score_0_x425;
      res_1_sum <= res_1_sum + score_1_x425;
      res_2_sum <= res_2_sum + score_2_x425;
      res_3_sum <= res_3_sum + score_3_x425;
      res_4_sum <= res_4_sum + score_4_x425;
      res_5_sum <= res_5_sum + score_5_x425;
      res_6_sum <= res_6_sum + score_6_x425;
      res_7_sum <= res_7_sum + score_7_x425;
      res_8_sum <= res_8_sum + score_8_x425;
      res_9_sum <= res_9_sum + score_9_x425;
   end
   else if(res_done_x426) begin
      res_0_sum <= res_0_sum + score_0_x426;
      res_1_sum <= res_1_sum + score_1_x426;
      res_2_sum <= res_2_sum + score_2_x426;
      res_3_sum <= res_3_sum + score_3_x426;
      res_4_sum <= res_4_sum + score_4_x426;
      res_5_sum <= res_5_sum + score_5_x426;
      res_6_sum <= res_6_sum + score_6_x426;
      res_7_sum <= res_7_sum + score_7_x426;
      res_8_sum <= res_8_sum + score_8_x426;
      res_9_sum <= res_9_sum + score_9_x426;
   end
   else if(res_done_x427) begin
      res_0_sum <= res_0_sum + score_0_x427;
      res_1_sum <= res_1_sum + score_1_x427;
      res_2_sum <= res_2_sum + score_2_x427;
      res_3_sum <= res_3_sum + score_3_x427;
      res_4_sum <= res_4_sum + score_4_x427;
      res_5_sum <= res_5_sum + score_5_x427;
      res_6_sum <= res_6_sum + score_6_x427;
      res_7_sum <= res_7_sum + score_7_x427;
      res_8_sum <= res_8_sum + score_8_x427;
      res_9_sum <= res_9_sum + score_9_x427;
   end
   else if(res_done_x428) begin
      res_0_sum <= res_0_sum + score_0_x428;
      res_1_sum <= res_1_sum + score_1_x428;
      res_2_sum <= res_2_sum + score_2_x428;
      res_3_sum <= res_3_sum + score_3_x428;
      res_4_sum <= res_4_sum + score_4_x428;
      res_5_sum <= res_5_sum + score_5_x428;
      res_6_sum <= res_6_sum + score_6_x428;
      res_7_sum <= res_7_sum + score_7_x428;
      res_8_sum <= res_8_sum + score_8_x428;
      res_9_sum <= res_9_sum + score_9_x428;
   end
   else if(res_done_x429) begin
      res_0_sum <= res_0_sum + score_0_x429;
      res_1_sum <= res_1_sum + score_1_x429;
      res_2_sum <= res_2_sum + score_2_x429;
      res_3_sum <= res_3_sum + score_3_x429;
      res_4_sum <= res_4_sum + score_4_x429;
      res_5_sum <= res_5_sum + score_5_x429;
      res_6_sum <= res_6_sum + score_6_x429;
      res_7_sum <= res_7_sum + score_7_x429;
      res_8_sum <= res_8_sum + score_8_x429;
      res_9_sum <= res_9_sum + score_9_x429;
   end
   else if(res_done_x430) begin
      res_0_sum <= res_0_sum + score_0_x430;
      res_1_sum <= res_1_sum + score_1_x430;
      res_2_sum <= res_2_sum + score_2_x430;
      res_3_sum <= res_3_sum + score_3_x430;
      res_4_sum <= res_4_sum + score_4_x430;
      res_5_sum <= res_5_sum + score_5_x430;
      res_6_sum <= res_6_sum + score_6_x430;
      res_7_sum <= res_7_sum + score_7_x430;
      res_8_sum <= res_8_sum + score_8_x430;
      res_9_sum <= res_9_sum + score_9_x430;
   end
   else if(res_done_x431) begin
      res_0_sum <= res_0_sum + score_0_x431;
      res_1_sum <= res_1_sum + score_1_x431;
      res_2_sum <= res_2_sum + score_2_x431;
      res_3_sum <= res_3_sum + score_3_x431;
      res_4_sum <= res_4_sum + score_4_x431;
      res_5_sum <= res_5_sum + score_5_x431;
      res_6_sum <= res_6_sum + score_6_x431;
      res_7_sum <= res_7_sum + score_7_x431;
      res_8_sum <= res_8_sum + score_8_x431;
      res_9_sum <= res_9_sum + score_9_x431;
   end
   else if(res_done_x432) begin
      res_0_sum <= res_0_sum + score_0_x432;
      res_1_sum <= res_1_sum + score_1_x432;
      res_2_sum <= res_2_sum + score_2_x432;
      res_3_sum <= res_3_sum + score_3_x432;
      res_4_sum <= res_4_sum + score_4_x432;
      res_5_sum <= res_5_sum + score_5_x432;
      res_6_sum <= res_6_sum + score_6_x432;
      res_7_sum <= res_7_sum + score_7_x432;
      res_8_sum <= res_8_sum + score_8_x432;
      res_9_sum <= res_9_sum + score_9_x432;
   end
   else if(res_done_x433) begin
      res_0_sum <= res_0_sum + score_0_x433;
      res_1_sum <= res_1_sum + score_1_x433;
      res_2_sum <= res_2_sum + score_2_x433;
      res_3_sum <= res_3_sum + score_3_x433;
      res_4_sum <= res_4_sum + score_4_x433;
      res_5_sum <= res_5_sum + score_5_x433;
      res_6_sum <= res_6_sum + score_6_x433;
      res_7_sum <= res_7_sum + score_7_x433;
      res_8_sum <= res_8_sum + score_8_x433;
      res_9_sum <= res_9_sum + score_9_x433;
   end
   else if(res_done_x434) begin
      res_0_sum <= res_0_sum + score_0_x434;
      res_1_sum <= res_1_sum + score_1_x434;
      res_2_sum <= res_2_sum + score_2_x434;
      res_3_sum <= res_3_sum + score_3_x434;
      res_4_sum <= res_4_sum + score_4_x434;
      res_5_sum <= res_5_sum + score_5_x434;
      res_6_sum <= res_6_sum + score_6_x434;
      res_7_sum <= res_7_sum + score_7_x434;
      res_8_sum <= res_8_sum + score_8_x434;
      res_9_sum <= res_9_sum + score_9_x434;
   end
   else if(res_done_x435) begin
      res_0_sum <= res_0_sum + score_0_x435;
      res_1_sum <= res_1_sum + score_1_x435;
      res_2_sum <= res_2_sum + score_2_x435;
      res_3_sum <= res_3_sum + score_3_x435;
      res_4_sum <= res_4_sum + score_4_x435;
      res_5_sum <= res_5_sum + score_5_x435;
      res_6_sum <= res_6_sum + score_6_x435;
      res_7_sum <= res_7_sum + score_7_x435;
      res_8_sum <= res_8_sum + score_8_x435;
      res_9_sum <= res_9_sum + score_9_x435;
   end
   else if(res_done_x436) begin
      res_0_sum <= res_0_sum + score_0_x436;
      res_1_sum <= res_1_sum + score_1_x436;
      res_2_sum <= res_2_sum + score_2_x436;
      res_3_sum <= res_3_sum + score_3_x436;
      res_4_sum <= res_4_sum + score_4_x436;
      res_5_sum <= res_5_sum + score_5_x436;
      res_6_sum <= res_6_sum + score_6_x436;
      res_7_sum <= res_7_sum + score_7_x436;
      res_8_sum <= res_8_sum + score_8_x436;
      res_9_sum <= res_9_sum + score_9_x436;
   end
   else if(res_done_x437) begin
      res_0_sum <= res_0_sum + score_0_x437;
      res_1_sum <= res_1_sum + score_1_x437;
      res_2_sum <= res_2_sum + score_2_x437;
      res_3_sum <= res_3_sum + score_3_x437;
      res_4_sum <= res_4_sum + score_4_x437;
      res_5_sum <= res_5_sum + score_5_x437;
      res_6_sum <= res_6_sum + score_6_x437;
      res_7_sum <= res_7_sum + score_7_x437;
      res_8_sum <= res_8_sum + score_8_x437;
      res_9_sum <= res_9_sum + score_9_x437;
   end
   else if(res_done_x438) begin
      res_0_sum <= res_0_sum + score_0_x438;
      res_1_sum <= res_1_sum + score_1_x438;
      res_2_sum <= res_2_sum + score_2_x438;
      res_3_sum <= res_3_sum + score_3_x438;
      res_4_sum <= res_4_sum + score_4_x438;
      res_5_sum <= res_5_sum + score_5_x438;
      res_6_sum <= res_6_sum + score_6_x438;
      res_7_sum <= res_7_sum + score_7_x438;
      res_8_sum <= res_8_sum + score_8_x438;
      res_9_sum <= res_9_sum + score_9_x438;
   end
   else if(res_done_x439) begin
      res_0_sum <= res_0_sum + score_0_x439;
      res_1_sum <= res_1_sum + score_1_x439;
      res_2_sum <= res_2_sum + score_2_x439;
      res_3_sum <= res_3_sum + score_3_x439;
      res_4_sum <= res_4_sum + score_4_x439;
      res_5_sum <= res_5_sum + score_5_x439;
      res_6_sum <= res_6_sum + score_6_x439;
      res_7_sum <= res_7_sum + score_7_x439;
      res_8_sum <= res_8_sum + score_8_x439;
      res_9_sum <= res_9_sum + score_9_x439;
   end
   else if(res_done_x440) begin
      res_0_sum <= res_0_sum + score_0_x440;
      res_1_sum <= res_1_sum + score_1_x440;
      res_2_sum <= res_2_sum + score_2_x440;
      res_3_sum <= res_3_sum + score_3_x440;
      res_4_sum <= res_4_sum + score_4_x440;
      res_5_sum <= res_5_sum + score_5_x440;
      res_6_sum <= res_6_sum + score_6_x440;
      res_7_sum <= res_7_sum + score_7_x440;
      res_8_sum <= res_8_sum + score_8_x440;
      res_9_sum <= res_9_sum + score_9_x440;
   end
   else if(res_done_x441) begin
      res_0_sum <= res_0_sum + score_0_x441;
      res_1_sum <= res_1_sum + score_1_x441;
      res_2_sum <= res_2_sum + score_2_x441;
      res_3_sum <= res_3_sum + score_3_x441;
      res_4_sum <= res_4_sum + score_4_x441;
      res_5_sum <= res_5_sum + score_5_x441;
      res_6_sum <= res_6_sum + score_6_x441;
      res_7_sum <= res_7_sum + score_7_x441;
      res_8_sum <= res_8_sum + score_8_x441;
      res_9_sum <= res_9_sum + score_9_x441;
   end
   else if(res_done_x442) begin
      res_0_sum <= res_0_sum + score_0_x442;
      res_1_sum <= res_1_sum + score_1_x442;
      res_2_sum <= res_2_sum + score_2_x442;
      res_3_sum <= res_3_sum + score_3_x442;
      res_4_sum <= res_4_sum + score_4_x442;
      res_5_sum <= res_5_sum + score_5_x442;
      res_6_sum <= res_6_sum + score_6_x442;
      res_7_sum <= res_7_sum + score_7_x442;
      res_8_sum <= res_8_sum + score_8_x442;
      res_9_sum <= res_9_sum + score_9_x442;
   end
   else if(res_done_x443) begin
      res_0_sum <= res_0_sum + score_0_x443;
      res_1_sum <= res_1_sum + score_1_x443;
      res_2_sum <= res_2_sum + score_2_x443;
      res_3_sum <= res_3_sum + score_3_x443;
      res_4_sum <= res_4_sum + score_4_x443;
      res_5_sum <= res_5_sum + score_5_x443;
      res_6_sum <= res_6_sum + score_6_x443;
      res_7_sum <= res_7_sum + score_7_x443;
      res_8_sum <= res_8_sum + score_8_x443;
      res_9_sum <= res_9_sum + score_9_x443;
   end
   else if(res_done_x444) begin
      res_0_sum <= res_0_sum + score_0_x444;
      res_1_sum <= res_1_sum + score_1_x444;
      res_2_sum <= res_2_sum + score_2_x444;
      res_3_sum <= res_3_sum + score_3_x444;
      res_4_sum <= res_4_sum + score_4_x444;
      res_5_sum <= res_5_sum + score_5_x444;
      res_6_sum <= res_6_sum + score_6_x444;
      res_7_sum <= res_7_sum + score_7_x444;
      res_8_sum <= res_8_sum + score_8_x444;
      res_9_sum <= res_9_sum + score_9_x444;
   end
   else if(res_done_x445) begin
      res_0_sum <= res_0_sum + score_0_x445;
      res_1_sum <= res_1_sum + score_1_x445;
      res_2_sum <= res_2_sum + score_2_x445;
      res_3_sum <= res_3_sum + score_3_x445;
      res_4_sum <= res_4_sum + score_4_x445;
      res_5_sum <= res_5_sum + score_5_x445;
      res_6_sum <= res_6_sum + score_6_x445;
      res_7_sum <= res_7_sum + score_7_x445;
      res_8_sum <= res_8_sum + score_8_x445;
      res_9_sum <= res_9_sum + score_9_x445;
   end
   else if(res_done_x446) begin
      res_0_sum <= res_0_sum + score_0_x446;
      res_1_sum <= res_1_sum + score_1_x446;
      res_2_sum <= res_2_sum + score_2_x446;
      res_3_sum <= res_3_sum + score_3_x446;
      res_4_sum <= res_4_sum + score_4_x446;
      res_5_sum <= res_5_sum + score_5_x446;
      res_6_sum <= res_6_sum + score_6_x446;
      res_7_sum <= res_7_sum + score_7_x446;
      res_8_sum <= res_8_sum + score_8_x446;
      res_9_sum <= res_9_sum + score_9_x446;
   end
   else if(res_done_x447) begin
      res_0_sum <= res_0_sum + score_0_x447;
      res_1_sum <= res_1_sum + score_1_x447;
      res_2_sum <= res_2_sum + score_2_x447;
      res_3_sum <= res_3_sum + score_3_x447;
      res_4_sum <= res_4_sum + score_4_x447;
      res_5_sum <= res_5_sum + score_5_x447;
      res_6_sum <= res_6_sum + score_6_x447;
      res_7_sum <= res_7_sum + score_7_x447;
      res_8_sum <= res_8_sum + score_8_x447;
      res_9_sum <= res_9_sum + score_9_x447;
   end
   else if(res_done_x448) begin
      res_0_sum <= res_0_sum + score_0_x448;
      res_1_sum <= res_1_sum + score_1_x448;
      res_2_sum <= res_2_sum + score_2_x448;
      res_3_sum <= res_3_sum + score_3_x448;
      res_4_sum <= res_4_sum + score_4_x448;
      res_5_sum <= res_5_sum + score_5_x448;
      res_6_sum <= res_6_sum + score_6_x448;
      res_7_sum <= res_7_sum + score_7_x448;
      res_8_sum <= res_8_sum + score_8_x448;
      res_9_sum <= res_9_sum + score_9_x448;
   end
   else if(res_done_x449) begin
      res_0_sum <= res_0_sum + score_0_x449;
      res_1_sum <= res_1_sum + score_1_x449;
      res_2_sum <= res_2_sum + score_2_x449;
      res_3_sum <= res_3_sum + score_3_x449;
      res_4_sum <= res_4_sum + score_4_x449;
      res_5_sum <= res_5_sum + score_5_x449;
      res_6_sum <= res_6_sum + score_6_x449;
      res_7_sum <= res_7_sum + score_7_x449;
      res_8_sum <= res_8_sum + score_8_x449;
      res_9_sum <= res_9_sum + score_9_x449;
   end
   else if(res_done_x450) begin
      res_0_sum <= res_0_sum + score_0_x450;
      res_1_sum <= res_1_sum + score_1_x450;
      res_2_sum <= res_2_sum + score_2_x450;
      res_3_sum <= res_3_sum + score_3_x450;
      res_4_sum <= res_4_sum + score_4_x450;
      res_5_sum <= res_5_sum + score_5_x450;
      res_6_sum <= res_6_sum + score_6_x450;
      res_7_sum <= res_7_sum + score_7_x450;
      res_8_sum <= res_8_sum + score_8_x450;
      res_9_sum <= res_9_sum + score_9_x450;
   end
   else if(res_done_x451) begin
      res_0_sum <= res_0_sum + score_0_x451;
      res_1_sum <= res_1_sum + score_1_x451;
      res_2_sum <= res_2_sum + score_2_x451;
      res_3_sum <= res_3_sum + score_3_x451;
      res_4_sum <= res_4_sum + score_4_x451;
      res_5_sum <= res_5_sum + score_5_x451;
      res_6_sum <= res_6_sum + score_6_x451;
      res_7_sum <= res_7_sum + score_7_x451;
      res_8_sum <= res_8_sum + score_8_x451;
      res_9_sum <= res_9_sum + score_9_x451;
   end
   else if(res_done_x452) begin
      res_0_sum <= res_0_sum + score_0_x452;
      res_1_sum <= res_1_sum + score_1_x452;
      res_2_sum <= res_2_sum + score_2_x452;
      res_3_sum <= res_3_sum + score_3_x452;
      res_4_sum <= res_4_sum + score_4_x452;
      res_5_sum <= res_5_sum + score_5_x452;
      res_6_sum <= res_6_sum + score_6_x452;
      res_7_sum <= res_7_sum + score_7_x452;
      res_8_sum <= res_8_sum + score_8_x452;
      res_9_sum <= res_9_sum + score_9_x452;
   end
   else if(res_done_x453) begin
      res_0_sum <= res_0_sum + score_0_x453;
      res_1_sum <= res_1_sum + score_1_x453;
      res_2_sum <= res_2_sum + score_2_x453;
      res_3_sum <= res_3_sum + score_3_x453;
      res_4_sum <= res_4_sum + score_4_x453;
      res_5_sum <= res_5_sum + score_5_x453;
      res_6_sum <= res_6_sum + score_6_x453;
      res_7_sum <= res_7_sum + score_7_x453;
      res_8_sum <= res_8_sum + score_8_x453;
      res_9_sum <= res_9_sum + score_9_x453;
   end
   else if(res_done_x454) begin
      res_0_sum <= res_0_sum + score_0_x454;
      res_1_sum <= res_1_sum + score_1_x454;
      res_2_sum <= res_2_sum + score_2_x454;
      res_3_sum <= res_3_sum + score_3_x454;
      res_4_sum <= res_4_sum + score_4_x454;
      res_5_sum <= res_5_sum + score_5_x454;
      res_6_sum <= res_6_sum + score_6_x454;
      res_7_sum <= res_7_sum + score_7_x454;
      res_8_sum <= res_8_sum + score_8_x454;
      res_9_sum <= res_9_sum + score_9_x454;
   end
   else if(res_done_x455) begin
      res_0_sum <= res_0_sum + score_0_x455;
      res_1_sum <= res_1_sum + score_1_x455;
      res_2_sum <= res_2_sum + score_2_x455;
      res_3_sum <= res_3_sum + score_3_x455;
      res_4_sum <= res_4_sum + score_4_x455;
      res_5_sum <= res_5_sum + score_5_x455;
      res_6_sum <= res_6_sum + score_6_x455;
      res_7_sum <= res_7_sum + score_7_x455;
      res_8_sum <= res_8_sum + score_8_x455;
      res_9_sum <= res_9_sum + score_9_x455;
   end
   else if(res_done_x456) begin
      res_0_sum <= res_0_sum + score_0_x456;
      res_1_sum <= res_1_sum + score_1_x456;
      res_2_sum <= res_2_sum + score_2_x456;
      res_3_sum <= res_3_sum + score_3_x456;
      res_4_sum <= res_4_sum + score_4_x456;
      res_5_sum <= res_5_sum + score_5_x456;
      res_6_sum <= res_6_sum + score_6_x456;
      res_7_sum <= res_7_sum + score_7_x456;
      res_8_sum <= res_8_sum + score_8_x456;
      res_9_sum <= res_9_sum + score_9_x456;
   end
   else if(res_done_x457) begin
      res_0_sum <= res_0_sum + score_0_x457;
      res_1_sum <= res_1_sum + score_1_x457;
      res_2_sum <= res_2_sum + score_2_x457;
      res_3_sum <= res_3_sum + score_3_x457;
      res_4_sum <= res_4_sum + score_4_x457;
      res_5_sum <= res_5_sum + score_5_x457;
      res_6_sum <= res_6_sum + score_6_x457;
      res_7_sum <= res_7_sum + score_7_x457;
      res_8_sum <= res_8_sum + score_8_x457;
      res_9_sum <= res_9_sum + score_9_x457;
   end
   else if(res_done_x458) begin
      res_0_sum <= res_0_sum + score_0_x458;
      res_1_sum <= res_1_sum + score_1_x458;
      res_2_sum <= res_2_sum + score_2_x458;
      res_3_sum <= res_3_sum + score_3_x458;
      res_4_sum <= res_4_sum + score_4_x458;
      res_5_sum <= res_5_sum + score_5_x458;
      res_6_sum <= res_6_sum + score_6_x458;
      res_7_sum <= res_7_sum + score_7_x458;
      res_8_sum <= res_8_sum + score_8_x458;
      res_9_sum <= res_9_sum + score_9_x458;
   end
   else if(res_done_x459) begin
      res_0_sum <= res_0_sum + score_0_x459;
      res_1_sum <= res_1_sum + score_1_x459;
      res_2_sum <= res_2_sum + score_2_x459;
      res_3_sum <= res_3_sum + score_3_x459;
      res_4_sum <= res_4_sum + score_4_x459;
      res_5_sum <= res_5_sum + score_5_x459;
      res_6_sum <= res_6_sum + score_6_x459;
      res_7_sum <= res_7_sum + score_7_x459;
      res_8_sum <= res_8_sum + score_8_x459;
      res_9_sum <= res_9_sum + score_9_x459;
   end
   else if(res_done_x460) begin
      res_0_sum <= res_0_sum + score_0_x460;
      res_1_sum <= res_1_sum + score_1_x460;
      res_2_sum <= res_2_sum + score_2_x460;
      res_3_sum <= res_3_sum + score_3_x460;
      res_4_sum <= res_4_sum + score_4_x460;
      res_5_sum <= res_5_sum + score_5_x460;
      res_6_sum <= res_6_sum + score_6_x460;
      res_7_sum <= res_7_sum + score_7_x460;
      res_8_sum <= res_8_sum + score_8_x460;
      res_9_sum <= res_9_sum + score_9_x460;
   end
   else if(res_done_x461) begin
      res_0_sum <= res_0_sum + score_0_x461;
      res_1_sum <= res_1_sum + score_1_x461;
      res_2_sum <= res_2_sum + score_2_x461;
      res_3_sum <= res_3_sum + score_3_x461;
      res_4_sum <= res_4_sum + score_4_x461;
      res_5_sum <= res_5_sum + score_5_x461;
      res_6_sum <= res_6_sum + score_6_x461;
      res_7_sum <= res_7_sum + score_7_x461;
      res_8_sum <= res_8_sum + score_8_x461;
      res_9_sum <= res_9_sum + score_9_x461;
   end
   else if(res_done_x462) begin
      res_0_sum <= res_0_sum + score_0_x462;
      res_1_sum <= res_1_sum + score_1_x462;
      res_2_sum <= res_2_sum + score_2_x462;
      res_3_sum <= res_3_sum + score_3_x462;
      res_4_sum <= res_4_sum + score_4_x462;
      res_5_sum <= res_5_sum + score_5_x462;
      res_6_sum <= res_6_sum + score_6_x462;
      res_7_sum <= res_7_sum + score_7_x462;
      res_8_sum <= res_8_sum + score_8_x462;
      res_9_sum <= res_9_sum + score_9_x462;
   end
   else if(res_done_x463) begin
      res_0_sum <= res_0_sum + score_0_x463;
      res_1_sum <= res_1_sum + score_1_x463;
      res_2_sum <= res_2_sum + score_2_x463;
      res_3_sum <= res_3_sum + score_3_x463;
      res_4_sum <= res_4_sum + score_4_x463;
      res_5_sum <= res_5_sum + score_5_x463;
      res_6_sum <= res_6_sum + score_6_x463;
      res_7_sum <= res_7_sum + score_7_x463;
      res_8_sum <= res_8_sum + score_8_x463;
      res_9_sum <= res_9_sum + score_9_x463;
   end
   else if(res_done_x464) begin
      res_0_sum <= res_0_sum + score_0_x464;
      res_1_sum <= res_1_sum + score_1_x464;
      res_2_sum <= res_2_sum + score_2_x464;
      res_3_sum <= res_3_sum + score_3_x464;
      res_4_sum <= res_4_sum + score_4_x464;
      res_5_sum <= res_5_sum + score_5_x464;
      res_6_sum <= res_6_sum + score_6_x464;
      res_7_sum <= res_7_sum + score_7_x464;
      res_8_sum <= res_8_sum + score_8_x464;
      res_9_sum <= res_9_sum + score_9_x464;
   end
   else if(res_done_x465) begin
      res_0_sum <= res_0_sum + score_0_x465;
      res_1_sum <= res_1_sum + score_1_x465;
      res_2_sum <= res_2_sum + score_2_x465;
      res_3_sum <= res_3_sum + score_3_x465;
      res_4_sum <= res_4_sum + score_4_x465;
      res_5_sum <= res_5_sum + score_5_x465;
      res_6_sum <= res_6_sum + score_6_x465;
      res_7_sum <= res_7_sum + score_7_x465;
      res_8_sum <= res_8_sum + score_8_x465;
      res_9_sum <= res_9_sum + score_9_x465;
   end
   else if(res_done_x466) begin
      res_0_sum <= res_0_sum + score_0_x466;
      res_1_sum <= res_1_sum + score_1_x466;
      res_2_sum <= res_2_sum + score_2_x466;
      res_3_sum <= res_3_sum + score_3_x466;
      res_4_sum <= res_4_sum + score_4_x466;
      res_5_sum <= res_5_sum + score_5_x466;
      res_6_sum <= res_6_sum + score_6_x466;
      res_7_sum <= res_7_sum + score_7_x466;
      res_8_sum <= res_8_sum + score_8_x466;
      res_9_sum <= res_9_sum + score_9_x466;
   end
   else if(res_done_x467) begin
      res_0_sum <= res_0_sum + score_0_x467;
      res_1_sum <= res_1_sum + score_1_x467;
      res_2_sum <= res_2_sum + score_2_x467;
      res_3_sum <= res_3_sum + score_3_x467;
      res_4_sum <= res_4_sum + score_4_x467;
      res_5_sum <= res_5_sum + score_5_x467;
      res_6_sum <= res_6_sum + score_6_x467;
      res_7_sum <= res_7_sum + score_7_x467;
      res_8_sum <= res_8_sum + score_8_x467;
      res_9_sum <= res_9_sum + score_9_x467;
   end
   else if(res_done_x468) begin
      res_0_sum <= res_0_sum + score_0_x468;
      res_1_sum <= res_1_sum + score_1_x468;
      res_2_sum <= res_2_sum + score_2_x468;
      res_3_sum <= res_3_sum + score_3_x468;
      res_4_sum <= res_4_sum + score_4_x468;
      res_5_sum <= res_5_sum + score_5_x468;
      res_6_sum <= res_6_sum + score_6_x468;
      res_7_sum <= res_7_sum + score_7_x468;
      res_8_sum <= res_8_sum + score_8_x468;
      res_9_sum <= res_9_sum + score_9_x468;
   end
   else if(res_done_x469) begin
      res_0_sum <= res_0_sum + score_0_x469;
      res_1_sum <= res_1_sum + score_1_x469;
      res_2_sum <= res_2_sum + score_2_x469;
      res_3_sum <= res_3_sum + score_3_x469;
      res_4_sum <= res_4_sum + score_4_x469;
      res_5_sum <= res_5_sum + score_5_x469;
      res_6_sum <= res_6_sum + score_6_x469;
      res_7_sum <= res_7_sum + score_7_x469;
      res_8_sum <= res_8_sum + score_8_x469;
      res_9_sum <= res_9_sum + score_9_x469;
   end
   else if(res_done_x470) begin
      res_0_sum <= res_0_sum + score_0_x470;
      res_1_sum <= res_1_sum + score_1_x470;
      res_2_sum <= res_2_sum + score_2_x470;
      res_3_sum <= res_3_sum + score_3_x470;
      res_4_sum <= res_4_sum + score_4_x470;
      res_5_sum <= res_5_sum + score_5_x470;
      res_6_sum <= res_6_sum + score_6_x470;
      res_7_sum <= res_7_sum + score_7_x470;
      res_8_sum <= res_8_sum + score_8_x470;
      res_9_sum <= res_9_sum + score_9_x470;
   end
   else if(res_done_x471) begin
      res_0_sum <= res_0_sum + score_0_x471;
      res_1_sum <= res_1_sum + score_1_x471;
      res_2_sum <= res_2_sum + score_2_x471;
      res_3_sum <= res_3_sum + score_3_x471;
      res_4_sum <= res_4_sum + score_4_x471;
      res_5_sum <= res_5_sum + score_5_x471;
      res_6_sum <= res_6_sum + score_6_x471;
      res_7_sum <= res_7_sum + score_7_x471;
      res_8_sum <= res_8_sum + score_8_x471;
      res_9_sum <= res_9_sum + score_9_x471;
   end
   else if(res_done_x472) begin
      res_0_sum <= res_0_sum + score_0_x472;
      res_1_sum <= res_1_sum + score_1_x472;
      res_2_sum <= res_2_sum + score_2_x472;
      res_3_sum <= res_3_sum + score_3_x472;
      res_4_sum <= res_4_sum + score_4_x472;
      res_5_sum <= res_5_sum + score_5_x472;
      res_6_sum <= res_6_sum + score_6_x472;
      res_7_sum <= res_7_sum + score_7_x472;
      res_8_sum <= res_8_sum + score_8_x472;
      res_9_sum <= res_9_sum + score_9_x472;
   end
   else if(res_done_x473) begin
      res_0_sum <= res_0_sum + score_0_x473;
      res_1_sum <= res_1_sum + score_1_x473;
      res_2_sum <= res_2_sum + score_2_x473;
      res_3_sum <= res_3_sum + score_3_x473;
      res_4_sum <= res_4_sum + score_4_x473;
      res_5_sum <= res_5_sum + score_5_x473;
      res_6_sum <= res_6_sum + score_6_x473;
      res_7_sum <= res_7_sum + score_7_x473;
      res_8_sum <= res_8_sum + score_8_x473;
      res_9_sum <= res_9_sum + score_9_x473;
   end
   else if(res_done_x474) begin
      res_0_sum <= res_0_sum + score_0_x474;
      res_1_sum <= res_1_sum + score_1_x474;
      res_2_sum <= res_2_sum + score_2_x474;
      res_3_sum <= res_3_sum + score_3_x474;
      res_4_sum <= res_4_sum + score_4_x474;
      res_5_sum <= res_5_sum + score_5_x474;
      res_6_sum <= res_6_sum + score_6_x474;
      res_7_sum <= res_7_sum + score_7_x474;
      res_8_sum <= res_8_sum + score_8_x474;
      res_9_sum <= res_9_sum + score_9_x474;
   end
   else if(res_done_x475) begin
      res_0_sum <= res_0_sum + score_0_x475;
      res_1_sum <= res_1_sum + score_1_x475;
      res_2_sum <= res_2_sum + score_2_x475;
      res_3_sum <= res_3_sum + score_3_x475;
      res_4_sum <= res_4_sum + score_4_x475;
      res_5_sum <= res_5_sum + score_5_x475;
      res_6_sum <= res_6_sum + score_6_x475;
      res_7_sum <= res_7_sum + score_7_x475;
      res_8_sum <= res_8_sum + score_8_x475;
      res_9_sum <= res_9_sum + score_9_x475;
   end
   else if(res_done_x476) begin
      res_0_sum <= res_0_sum + score_0_x476;
      res_1_sum <= res_1_sum + score_1_x476;
      res_2_sum <= res_2_sum + score_2_x476;
      res_3_sum <= res_3_sum + score_3_x476;
      res_4_sum <= res_4_sum + score_4_x476;
      res_5_sum <= res_5_sum + score_5_x476;
      res_6_sum <= res_6_sum + score_6_x476;
      res_7_sum <= res_7_sum + score_7_x476;
      res_8_sum <= res_8_sum + score_8_x476;
      res_9_sum <= res_9_sum + score_9_x476;
   end
   else if(res_done_x477) begin
      res_0_sum <= res_0_sum + score_0_x477;
      res_1_sum <= res_1_sum + score_1_x477;
      res_2_sum <= res_2_sum + score_2_x477;
      res_3_sum <= res_3_sum + score_3_x477;
      res_4_sum <= res_4_sum + score_4_x477;
      res_5_sum <= res_5_sum + score_5_x477;
      res_6_sum <= res_6_sum + score_6_x477;
      res_7_sum <= res_7_sum + score_7_x477;
      res_8_sum <= res_8_sum + score_8_x477;
      res_9_sum <= res_9_sum + score_9_x477;
   end
   else if(res_done_x478) begin
      res_0_sum <= res_0_sum + score_0_x478;
      res_1_sum <= res_1_sum + score_1_x478;
      res_2_sum <= res_2_sum + score_2_x478;
      res_3_sum <= res_3_sum + score_3_x478;
      res_4_sum <= res_4_sum + score_4_x478;
      res_5_sum <= res_5_sum + score_5_x478;
      res_6_sum <= res_6_sum + score_6_x478;
      res_7_sum <= res_7_sum + score_7_x478;
      res_8_sum <= res_8_sum + score_8_x478;
      res_9_sum <= res_9_sum + score_9_x478;
   end
   else if(res_done_x479) begin
      res_0_sum <= res_0_sum + score_0_x479;
      res_1_sum <= res_1_sum + score_1_x479;
      res_2_sum <= res_2_sum + score_2_x479;
      res_3_sum <= res_3_sum + score_3_x479;
      res_4_sum <= res_4_sum + score_4_x479;
      res_5_sum <= res_5_sum + score_5_x479;
      res_6_sum <= res_6_sum + score_6_x479;
      res_7_sum <= res_7_sum + score_7_x479;
      res_8_sum <= res_8_sum + score_8_x479;
      res_9_sum <= res_9_sum + score_9_x479;
   end
   else if(res_done_x480) begin
      res_0_sum <= res_0_sum + score_0_x480;
      res_1_sum <= res_1_sum + score_1_x480;
      res_2_sum <= res_2_sum + score_2_x480;
      res_3_sum <= res_3_sum + score_3_x480;
      res_4_sum <= res_4_sum + score_4_x480;
      res_5_sum <= res_5_sum + score_5_x480;
      res_6_sum <= res_6_sum + score_6_x480;
      res_7_sum <= res_7_sum + score_7_x480;
      res_8_sum <= res_8_sum + score_8_x480;
      res_9_sum <= res_9_sum + score_9_x480;
   end
   else if(res_done_x481) begin
      res_0_sum <= res_0_sum + score_0_x481;
      res_1_sum <= res_1_sum + score_1_x481;
      res_2_sum <= res_2_sum + score_2_x481;
      res_3_sum <= res_3_sum + score_3_x481;
      res_4_sum <= res_4_sum + score_4_x481;
      res_5_sum <= res_5_sum + score_5_x481;
      res_6_sum <= res_6_sum + score_6_x481;
      res_7_sum <= res_7_sum + score_7_x481;
      res_8_sum <= res_8_sum + score_8_x481;
      res_9_sum <= res_9_sum + score_9_x481;
   end
   else if(res_done_x482) begin
      res_0_sum <= res_0_sum + score_0_x482;
      res_1_sum <= res_1_sum + score_1_x482;
      res_2_sum <= res_2_sum + score_2_x482;
      res_3_sum <= res_3_sum + score_3_x482;
      res_4_sum <= res_4_sum + score_4_x482;
      res_5_sum <= res_5_sum + score_5_x482;
      res_6_sum <= res_6_sum + score_6_x482;
      res_7_sum <= res_7_sum + score_7_x482;
      res_8_sum <= res_8_sum + score_8_x482;
      res_9_sum <= res_9_sum + score_9_x482;
   end
   else if(res_done_x483) begin
      res_0_sum <= res_0_sum + score_0_x483;
      res_1_sum <= res_1_sum + score_1_x483;
      res_2_sum <= res_2_sum + score_2_x483;
      res_3_sum <= res_3_sum + score_3_x483;
      res_4_sum <= res_4_sum + score_4_x483;
      res_5_sum <= res_5_sum + score_5_x483;
      res_6_sum <= res_6_sum + score_6_x483;
      res_7_sum <= res_7_sum + score_7_x483;
      res_8_sum <= res_8_sum + score_8_x483;
      res_9_sum <= res_9_sum + score_9_x483;
   end
   else if(res_done_x484) begin
      res_0_sum <= res_0_sum + score_0_x484;
      res_1_sum <= res_1_sum + score_1_x484;
      res_2_sum <= res_2_sum + score_2_x484;
      res_3_sum <= res_3_sum + score_3_x484;
      res_4_sum <= res_4_sum + score_4_x484;
      res_5_sum <= res_5_sum + score_5_x484;
      res_6_sum <= res_6_sum + score_6_x484;
      res_7_sum <= res_7_sum + score_7_x484;
      res_8_sum <= res_8_sum + score_8_x484;
      res_9_sum <= res_9_sum + score_9_x484;
   end
   else if(res_done_x485) begin
      res_0_sum <= res_0_sum + score_0_x485;
      res_1_sum <= res_1_sum + score_1_x485;
      res_2_sum <= res_2_sum + score_2_x485;
      res_3_sum <= res_3_sum + score_3_x485;
      res_4_sum <= res_4_sum + score_4_x485;
      res_5_sum <= res_5_sum + score_5_x485;
      res_6_sum <= res_6_sum + score_6_x485;
      res_7_sum <= res_7_sum + score_7_x485;
      res_8_sum <= res_8_sum + score_8_x485;
      res_9_sum <= res_9_sum + score_9_x485;
   end
   else if(res_done_x486) begin
      res_0_sum <= res_0_sum + score_0_x486;
      res_1_sum <= res_1_sum + score_1_x486;
      res_2_sum <= res_2_sum + score_2_x486;
      res_3_sum <= res_3_sum + score_3_x486;
      res_4_sum <= res_4_sum + score_4_x486;
      res_5_sum <= res_5_sum + score_5_x486;
      res_6_sum <= res_6_sum + score_6_x486;
      res_7_sum <= res_7_sum + score_7_x486;
      res_8_sum <= res_8_sum + score_8_x486;
      res_9_sum <= res_9_sum + score_9_x486;
   end
   else if(res_done_x487) begin
      res_0_sum <= res_0_sum + score_0_x487;
      res_1_sum <= res_1_sum + score_1_x487;
      res_2_sum <= res_2_sum + score_2_x487;
      res_3_sum <= res_3_sum + score_3_x487;
      res_4_sum <= res_4_sum + score_4_x487;
      res_5_sum <= res_5_sum + score_5_x487;
      res_6_sum <= res_6_sum + score_6_x487;
      res_7_sum <= res_7_sum + score_7_x487;
      res_8_sum <= res_8_sum + score_8_x487;
      res_9_sum <= res_9_sum + score_9_x487;
   end
   else if(res_done_x488) begin
      res_0_sum <= res_0_sum + score_0_x488;
      res_1_sum <= res_1_sum + score_1_x488;
      res_2_sum <= res_2_sum + score_2_x488;
      res_3_sum <= res_3_sum + score_3_x488;
      res_4_sum <= res_4_sum + score_4_x488;
      res_5_sum <= res_5_sum + score_5_x488;
      res_6_sum <= res_6_sum + score_6_x488;
      res_7_sum <= res_7_sum + score_7_x488;
      res_8_sum <= res_8_sum + score_8_x488;
      res_9_sum <= res_9_sum + score_9_x488;
   end
   else if(res_done_x489) begin
      res_0_sum <= res_0_sum + score_0_x489;
      res_1_sum <= res_1_sum + score_1_x489;
      res_2_sum <= res_2_sum + score_2_x489;
      res_3_sum <= res_3_sum + score_3_x489;
      res_4_sum <= res_4_sum + score_4_x489;
      res_5_sum <= res_5_sum + score_5_x489;
      res_6_sum <= res_6_sum + score_6_x489;
      res_7_sum <= res_7_sum + score_7_x489;
      res_8_sum <= res_8_sum + score_8_x489;
      res_9_sum <= res_9_sum + score_9_x489;
   end
   else if(res_done_x490) begin
      res_0_sum <= res_0_sum + score_0_x490;
      res_1_sum <= res_1_sum + score_1_x490;
      res_2_sum <= res_2_sum + score_2_x490;
      res_3_sum <= res_3_sum + score_3_x490;
      res_4_sum <= res_4_sum + score_4_x490;
      res_5_sum <= res_5_sum + score_5_x490;
      res_6_sum <= res_6_sum + score_6_x490;
      res_7_sum <= res_7_sum + score_7_x490;
      res_8_sum <= res_8_sum + score_8_x490;
      res_9_sum <= res_9_sum + score_9_x490;
   end
   else if(res_done_x491) begin
      res_0_sum <= res_0_sum + score_0_x491;
      res_1_sum <= res_1_sum + score_1_x491;
      res_2_sum <= res_2_sum + score_2_x491;
      res_3_sum <= res_3_sum + score_3_x491;
      res_4_sum <= res_4_sum + score_4_x491;
      res_5_sum <= res_5_sum + score_5_x491;
      res_6_sum <= res_6_sum + score_6_x491;
      res_7_sum <= res_7_sum + score_7_x491;
      res_8_sum <= res_8_sum + score_8_x491;
      res_9_sum <= res_9_sum + score_9_x491;
   end
   else if(res_done_x492) begin
      res_0_sum <= res_0_sum + score_0_x492;
      res_1_sum <= res_1_sum + score_1_x492;
      res_2_sum <= res_2_sum + score_2_x492;
      res_3_sum <= res_3_sum + score_3_x492;
      res_4_sum <= res_4_sum + score_4_x492;
      res_5_sum <= res_5_sum + score_5_x492;
      res_6_sum <= res_6_sum + score_6_x492;
      res_7_sum <= res_7_sum + score_7_x492;
      res_8_sum <= res_8_sum + score_8_x492;
      res_9_sum <= res_9_sum + score_9_x492;
   end
   else if(res_done_x493) begin
      res_0_sum <= res_0_sum + score_0_x493;
      res_1_sum <= res_1_sum + score_1_x493;
      res_2_sum <= res_2_sum + score_2_x493;
      res_3_sum <= res_3_sum + score_3_x493;
      res_4_sum <= res_4_sum + score_4_x493;
      res_5_sum <= res_5_sum + score_5_x493;
      res_6_sum <= res_6_sum + score_6_x493;
      res_7_sum <= res_7_sum + score_7_x493;
      res_8_sum <= res_8_sum + score_8_x493;
      res_9_sum <= res_9_sum + score_9_x493;
   end
   else if(res_done_x494) begin
      res_0_sum <= res_0_sum + score_0_x494;
      res_1_sum <= res_1_sum + score_1_x494;
      res_2_sum <= res_2_sum + score_2_x494;
      res_3_sum <= res_3_sum + score_3_x494;
      res_4_sum <= res_4_sum + score_4_x494;
      res_5_sum <= res_5_sum + score_5_x494;
      res_6_sum <= res_6_sum + score_6_x494;
      res_7_sum <= res_7_sum + score_7_x494;
      res_8_sum <= res_8_sum + score_8_x494;
      res_9_sum <= res_9_sum + score_9_x494;
   end
   else if(res_done_x495) begin
      res_0_sum <= res_0_sum + score_0_x495;
      res_1_sum <= res_1_sum + score_1_x495;
      res_2_sum <= res_2_sum + score_2_x495;
      res_3_sum <= res_3_sum + score_3_x495;
      res_4_sum <= res_4_sum + score_4_x495;
      res_5_sum <= res_5_sum + score_5_x495;
      res_6_sum <= res_6_sum + score_6_x495;
      res_7_sum <= res_7_sum + score_7_x495;
      res_8_sum <= res_8_sum + score_8_x495;
      res_9_sum <= res_9_sum + score_9_x495;
   end
   else if(res_done_x496) begin
      res_0_sum <= res_0_sum + score_0_x496;
      res_1_sum <= res_1_sum + score_1_x496;
      res_2_sum <= res_2_sum + score_2_x496;
      res_3_sum <= res_3_sum + score_3_x496;
      res_4_sum <= res_4_sum + score_4_x496;
      res_5_sum <= res_5_sum + score_5_x496;
      res_6_sum <= res_6_sum + score_6_x496;
      res_7_sum <= res_7_sum + score_7_x496;
      res_8_sum <= res_8_sum + score_8_x496;
      res_9_sum <= res_9_sum + score_9_x496;
   end
   else if(res_done_x497) begin
      res_0_sum <= res_0_sum + score_0_x497;
      res_1_sum <= res_1_sum + score_1_x497;
      res_2_sum <= res_2_sum + score_2_x497;
      res_3_sum <= res_3_sum + score_3_x497;
      res_4_sum <= res_4_sum + score_4_x497;
      res_5_sum <= res_5_sum + score_5_x497;
      res_6_sum <= res_6_sum + score_6_x497;
      res_7_sum <= res_7_sum + score_7_x497;
      res_8_sum <= res_8_sum + score_8_x497;
      res_9_sum <= res_9_sum + score_9_x497;
   end
   else if(res_done_x498) begin
      res_0_sum <= res_0_sum + score_0_x498;
      res_1_sum <= res_1_sum + score_1_x498;
      res_2_sum <= res_2_sum + score_2_x498;
      res_3_sum <= res_3_sum + score_3_x498;
      res_4_sum <= res_4_sum + score_4_x498;
      res_5_sum <= res_5_sum + score_5_x498;
      res_6_sum <= res_6_sum + score_6_x498;
      res_7_sum <= res_7_sum + score_7_x498;
      res_8_sum <= res_8_sum + score_8_x498;
      res_9_sum <= res_9_sum + score_9_x498;
   end
   else if(res_done_x499) begin
      res_0_sum <= res_0_sum + score_0_x499;
      res_1_sum <= res_1_sum + score_1_x499;
      res_2_sum <= res_2_sum + score_2_x499;
      res_3_sum <= res_3_sum + score_3_x499;
      res_4_sum <= res_4_sum + score_4_x499;
      res_5_sum <= res_5_sum + score_5_x499;
      res_6_sum <= res_6_sum + score_6_x499;
      res_7_sum <= res_7_sum + score_7_x499;
      res_8_sum <= res_8_sum + score_8_x499;
      res_9_sum <= res_9_sum + score_9_x499;
   end
   else if(res_done_x500) begin
      res_0_sum <= res_0_sum + score_0_x500;
      res_1_sum <= res_1_sum + score_1_x500;
      res_2_sum <= res_2_sum + score_2_x500;
      res_3_sum <= res_3_sum + score_3_x500;
      res_4_sum <= res_4_sum + score_4_x500;
      res_5_sum <= res_5_sum + score_5_x500;
      res_6_sum <= res_6_sum + score_6_x500;
      res_7_sum <= res_7_sum + score_7_x500;
      res_8_sum <= res_8_sum + score_8_x500;
      res_9_sum <= res_9_sum + score_9_x500;
   end
   else if(res_done_x501) begin
      res_0_sum <= res_0_sum + score_0_x501;
      res_1_sum <= res_1_sum + score_1_x501;
      res_2_sum <= res_2_sum + score_2_x501;
      res_3_sum <= res_3_sum + score_3_x501;
      res_4_sum <= res_4_sum + score_4_x501;
      res_5_sum <= res_5_sum + score_5_x501;
      res_6_sum <= res_6_sum + score_6_x501;
      res_7_sum <= res_7_sum + score_7_x501;
      res_8_sum <= res_8_sum + score_8_x501;
      res_9_sum <= res_9_sum + score_9_x501;
   end
   else if(res_done_x502) begin
      res_0_sum <= res_0_sum + score_0_x502;
      res_1_sum <= res_1_sum + score_1_x502;
      res_2_sum <= res_2_sum + score_2_x502;
      res_3_sum <= res_3_sum + score_3_x502;
      res_4_sum <= res_4_sum + score_4_x502;
      res_5_sum <= res_5_sum + score_5_x502;
      res_6_sum <= res_6_sum + score_6_x502;
      res_7_sum <= res_7_sum + score_7_x502;
      res_8_sum <= res_8_sum + score_8_x502;
      res_9_sum <= res_9_sum + score_9_x502;
   end
   else if(res_done_x503) begin
      res_0_sum <= res_0_sum + score_0_x503;
      res_1_sum <= res_1_sum + score_1_x503;
      res_2_sum <= res_2_sum + score_2_x503;
      res_3_sum <= res_3_sum + score_3_x503;
      res_4_sum <= res_4_sum + score_4_x503;
      res_5_sum <= res_5_sum + score_5_x503;
      res_6_sum <= res_6_sum + score_6_x503;
      res_7_sum <= res_7_sum + score_7_x503;
      res_8_sum <= res_8_sum + score_8_x503;
      res_9_sum <= res_9_sum + score_9_x503;
   end
   else if(res_done_x504) begin
      res_0_sum <= res_0_sum + score_0_x504;
      res_1_sum <= res_1_sum + score_1_x504;
      res_2_sum <= res_2_sum + score_2_x504;
      res_3_sum <= res_3_sum + score_3_x504;
      res_4_sum <= res_4_sum + score_4_x504;
      res_5_sum <= res_5_sum + score_5_x504;
      res_6_sum <= res_6_sum + score_6_x504;
      res_7_sum <= res_7_sum + score_7_x504;
      res_8_sum <= res_8_sum + score_8_x504;
      res_9_sum <= res_9_sum + score_9_x504;
   end
   else if(res_done_x505) begin
      res_0_sum <= res_0_sum + score_0_x505;
      res_1_sum <= res_1_sum + score_1_x505;
      res_2_sum <= res_2_sum + score_2_x505;
      res_3_sum <= res_3_sum + score_3_x505;
      res_4_sum <= res_4_sum + score_4_x505;
      res_5_sum <= res_5_sum + score_5_x505;
      res_6_sum <= res_6_sum + score_6_x505;
      res_7_sum <= res_7_sum + score_7_x505;
      res_8_sum <= res_8_sum + score_8_x505;
      res_9_sum <= res_9_sum + score_9_x505;
   end
   else if(res_done_x506) begin
      res_0_sum <= res_0_sum + score_0_x506;
      res_1_sum <= res_1_sum + score_1_x506;
      res_2_sum <= res_2_sum + score_2_x506;
      res_3_sum <= res_3_sum + score_3_x506;
      res_4_sum <= res_4_sum + score_4_x506;
      res_5_sum <= res_5_sum + score_5_x506;
      res_6_sum <= res_6_sum + score_6_x506;
      res_7_sum <= res_7_sum + score_7_x506;
      res_8_sum <= res_8_sum + score_8_x506;
      res_9_sum <= res_9_sum + score_9_x506;
   end
   else if(res_done_x507) begin
      res_0_sum <= res_0_sum + score_0_x507;
      res_1_sum <= res_1_sum + score_1_x507;
      res_2_sum <= res_2_sum + score_2_x507;
      res_3_sum <= res_3_sum + score_3_x507;
      res_4_sum <= res_4_sum + score_4_x507;
      res_5_sum <= res_5_sum + score_5_x507;
      res_6_sum <= res_6_sum + score_6_x507;
      res_7_sum <= res_7_sum + score_7_x507;
      res_8_sum <= res_8_sum + score_8_x507;
      res_9_sum <= res_9_sum + score_9_x507;
   end
   else if(res_done_x508) begin
      res_0_sum <= res_0_sum + score_0_x508;
      res_1_sum <= res_1_sum + score_1_x508;
      res_2_sum <= res_2_sum + score_2_x508;
      res_3_sum <= res_3_sum + score_3_x508;
      res_4_sum <= res_4_sum + score_4_x508;
      res_5_sum <= res_5_sum + score_5_x508;
      res_6_sum <= res_6_sum + score_6_x508;
      res_7_sum <= res_7_sum + score_7_x508;
      res_8_sum <= res_8_sum + score_8_x508;
      res_9_sum <= res_9_sum + score_9_x508;
   end
   else if(res_done_x509) begin
      res_0_sum <= res_0_sum + score_0_x509;
      res_1_sum <= res_1_sum + score_1_x509;
      res_2_sum <= res_2_sum + score_2_x509;
      res_3_sum <= res_3_sum + score_3_x509;
      res_4_sum <= res_4_sum + score_4_x509;
      res_5_sum <= res_5_sum + score_5_x509;
      res_6_sum <= res_6_sum + score_6_x509;
      res_7_sum <= res_7_sum + score_7_x509;
      res_8_sum <= res_8_sum + score_8_x509;
      res_9_sum <= res_9_sum + score_9_x509;
   end
   else if(res_done_x510) begin
      res_0_sum <= res_0_sum + score_0_x510;
      res_1_sum <= res_1_sum + score_1_x510;
      res_2_sum <= res_2_sum + score_2_x510;
      res_3_sum <= res_3_sum + score_3_x510;
      res_4_sum <= res_4_sum + score_4_x510;
      res_5_sum <= res_5_sum + score_5_x510;
      res_6_sum <= res_6_sum + score_6_x510;
      res_7_sum <= res_7_sum + score_7_x510;
      res_8_sum <= res_8_sum + score_8_x510;
      res_9_sum <= res_9_sum + score_9_x510;
   end
   else if(res_done_x511) begin
      res_0_sum <= res_0_sum + score_0_x511;
      res_1_sum <= res_1_sum + score_1_x511;
      res_2_sum <= res_2_sum + score_2_x511;
      res_3_sum <= res_3_sum + score_3_x511;
      res_4_sum <= res_4_sum + score_4_x511;
      res_5_sum <= res_5_sum + score_5_x511;
      res_6_sum <= res_6_sum + score_6_x511;
      res_7_sum <= res_7_sum + score_7_x511;
      res_8_sum <= res_8_sum + score_8_x511;
      res_9_sum <= res_9_sum + score_9_x511;
   end
   else if(res_done_x512) begin
      res_0_sum <= res_0_sum + score_0_x512;
      res_1_sum <= res_1_sum + score_1_x512;
      res_2_sum <= res_2_sum + score_2_x512;
      res_3_sum <= res_3_sum + score_3_x512;
      res_4_sum <= res_4_sum + score_4_x512;
      res_5_sum <= res_5_sum + score_5_x512;
      res_6_sum <= res_6_sum + score_6_x512;
      res_7_sum <= res_7_sum + score_7_x512;
      res_8_sum <= res_8_sum + score_8_x512;
      res_9_sum <= res_9_sum + score_9_x512;
   end
   else if(res_done_x513) begin
      res_0_sum <= res_0_sum + score_0_x513;
      res_1_sum <= res_1_sum + score_1_x513;
      res_2_sum <= res_2_sum + score_2_x513;
      res_3_sum <= res_3_sum + score_3_x513;
      res_4_sum <= res_4_sum + score_4_x513;
      res_5_sum <= res_5_sum + score_5_x513;
      res_6_sum <= res_6_sum + score_6_x513;
      res_7_sum <= res_7_sum + score_7_x513;
      res_8_sum <= res_8_sum + score_8_x513;
      res_9_sum <= res_9_sum + score_9_x513;
   end
   else if(res_done_x514) begin
      res_0_sum <= res_0_sum + score_0_x514;
      res_1_sum <= res_1_sum + score_1_x514;
      res_2_sum <= res_2_sum + score_2_x514;
      res_3_sum <= res_3_sum + score_3_x514;
      res_4_sum <= res_4_sum + score_4_x514;
      res_5_sum <= res_5_sum + score_5_x514;
      res_6_sum <= res_6_sum + score_6_x514;
      res_7_sum <= res_7_sum + score_7_x514;
      res_8_sum <= res_8_sum + score_8_x514;
      res_9_sum <= res_9_sum + score_9_x514;
   end
   else if(res_done_x515) begin
      res_0_sum <= res_0_sum + score_0_x515;
      res_1_sum <= res_1_sum + score_1_x515;
      res_2_sum <= res_2_sum + score_2_x515;
      res_3_sum <= res_3_sum + score_3_x515;
      res_4_sum <= res_4_sum + score_4_x515;
      res_5_sum <= res_5_sum + score_5_x515;
      res_6_sum <= res_6_sum + score_6_x515;
      res_7_sum <= res_7_sum + score_7_x515;
      res_8_sum <= res_8_sum + score_8_x515;
      res_9_sum <= res_9_sum + score_9_x515;
   end
   else if(res_done_x516) begin
      res_0_sum <= res_0_sum + score_0_x516;
      res_1_sum <= res_1_sum + score_1_x516;
      res_2_sum <= res_2_sum + score_2_x516;
      res_3_sum <= res_3_sum + score_3_x516;
      res_4_sum <= res_4_sum + score_4_x516;
      res_5_sum <= res_5_sum + score_5_x516;
      res_6_sum <= res_6_sum + score_6_x516;
      res_7_sum <= res_7_sum + score_7_x516;
      res_8_sum <= res_8_sum + score_8_x516;
      res_9_sum <= res_9_sum + score_9_x516;
   end
   else if(res_done_x517) begin
      res_0_sum <= res_0_sum + score_0_x517;
      res_1_sum <= res_1_sum + score_1_x517;
      res_2_sum <= res_2_sum + score_2_x517;
      res_3_sum <= res_3_sum + score_3_x517;
      res_4_sum <= res_4_sum + score_4_x517;
      res_5_sum <= res_5_sum + score_5_x517;
      res_6_sum <= res_6_sum + score_6_x517;
      res_7_sum <= res_7_sum + score_7_x517;
      res_8_sum <= res_8_sum + score_8_x517;
      res_9_sum <= res_9_sum + score_9_x517;
   end
   else if(res_done_x518) begin
      res_0_sum <= res_0_sum + score_0_x518;
      res_1_sum <= res_1_sum + score_1_x518;
      res_2_sum <= res_2_sum + score_2_x518;
      res_3_sum <= res_3_sum + score_3_x518;
      res_4_sum <= res_4_sum + score_4_x518;
      res_5_sum <= res_5_sum + score_5_x518;
      res_6_sum <= res_6_sum + score_6_x518;
      res_7_sum <= res_7_sum + score_7_x518;
      res_8_sum <= res_8_sum + score_8_x518;
      res_9_sum <= res_9_sum + score_9_x518;
   end
   else if(res_done_x519) begin
      res_0_sum <= res_0_sum + score_0_x519;
      res_1_sum <= res_1_sum + score_1_x519;
      res_2_sum <= res_2_sum + score_2_x519;
      res_3_sum <= res_3_sum + score_3_x519;
      res_4_sum <= res_4_sum + score_4_x519;
      res_5_sum <= res_5_sum + score_5_x519;
      res_6_sum <= res_6_sum + score_6_x519;
      res_7_sum <= res_7_sum + score_7_x519;
      res_8_sum <= res_8_sum + score_8_x519;
      res_9_sum <= res_9_sum + score_9_x519;
   end
   else if(res_done_x520) begin
      res_0_sum <= res_0_sum + score_0_x520;
      res_1_sum <= res_1_sum + score_1_x520;
      res_2_sum <= res_2_sum + score_2_x520;
      res_3_sum <= res_3_sum + score_3_x520;
      res_4_sum <= res_4_sum + score_4_x520;
      res_5_sum <= res_5_sum + score_5_x520;
      res_6_sum <= res_6_sum + score_6_x520;
      res_7_sum <= res_7_sum + score_7_x520;
      res_8_sum <= res_8_sum + score_8_x520;
      res_9_sum <= res_9_sum + score_9_x520;
   end
   else if(res_done_x521) begin
      res_0_sum <= res_0_sum + score_0_x521;
      res_1_sum <= res_1_sum + score_1_x521;
      res_2_sum <= res_2_sum + score_2_x521;
      res_3_sum <= res_3_sum + score_3_x521;
      res_4_sum <= res_4_sum + score_4_x521;
      res_5_sum <= res_5_sum + score_5_x521;
      res_6_sum <= res_6_sum + score_6_x521;
      res_7_sum <= res_7_sum + score_7_x521;
      res_8_sum <= res_8_sum + score_8_x521;
      res_9_sum <= res_9_sum + score_9_x521;
   end
   else if(res_done_x522) begin
      res_0_sum <= res_0_sum + score_0_x522;
      res_1_sum <= res_1_sum + score_1_x522;
      res_2_sum <= res_2_sum + score_2_x522;
      res_3_sum <= res_3_sum + score_3_x522;
      res_4_sum <= res_4_sum + score_4_x522;
      res_5_sum <= res_5_sum + score_5_x522;
      res_6_sum <= res_6_sum + score_6_x522;
      res_7_sum <= res_7_sum + score_7_x522;
      res_8_sum <= res_8_sum + score_8_x522;
      res_9_sum <= res_9_sum + score_9_x522;
   end
   else if(res_done_x523) begin
      res_0_sum <= res_0_sum + score_0_x523;
      res_1_sum <= res_1_sum + score_1_x523;
      res_2_sum <= res_2_sum + score_2_x523;
      res_3_sum <= res_3_sum + score_3_x523;
      res_4_sum <= res_4_sum + score_4_x523;
      res_5_sum <= res_5_sum + score_5_x523;
      res_6_sum <= res_6_sum + score_6_x523;
      res_7_sum <= res_7_sum + score_7_x523;
      res_8_sum <= res_8_sum + score_8_x523;
      res_9_sum <= res_9_sum + score_9_x523;
   end
   else if(res_done_x524) begin
      res_0_sum <= res_0_sum + score_0_x524;
      res_1_sum <= res_1_sum + score_1_x524;
      res_2_sum <= res_2_sum + score_2_x524;
      res_3_sum <= res_3_sum + score_3_x524;
      res_4_sum <= res_4_sum + score_4_x524;
      res_5_sum <= res_5_sum + score_5_x524;
      res_6_sum <= res_6_sum + score_6_x524;
      res_7_sum <= res_7_sum + score_7_x524;
      res_8_sum <= res_8_sum + score_8_x524;
      res_9_sum <= res_9_sum + score_9_x524;
   end
   else if(res_done_x525) begin
      res_0_sum <= res_0_sum + score_0_x525;
      res_1_sum <= res_1_sum + score_1_x525;
      res_2_sum <= res_2_sum + score_2_x525;
      res_3_sum <= res_3_sum + score_3_x525;
      res_4_sum <= res_4_sum + score_4_x525;
      res_5_sum <= res_5_sum + score_5_x525;
      res_6_sum <= res_6_sum + score_6_x525;
      res_7_sum <= res_7_sum + score_7_x525;
      res_8_sum <= res_8_sum + score_8_x525;
      res_9_sum <= res_9_sum + score_9_x525;
   end
   else if(res_done_x526) begin
      res_0_sum <= res_0_sum + score_0_x526;
      res_1_sum <= res_1_sum + score_1_x526;
      res_2_sum <= res_2_sum + score_2_x526;
      res_3_sum <= res_3_sum + score_3_x526;
      res_4_sum <= res_4_sum + score_4_x526;
      res_5_sum <= res_5_sum + score_5_x526;
      res_6_sum <= res_6_sum + score_6_x526;
      res_7_sum <= res_7_sum + score_7_x526;
      res_8_sum <= res_8_sum + score_8_x526;
      res_9_sum <= res_9_sum + score_9_x526;
   end
   else if(res_done_x527) begin
      res_0_sum <= res_0_sum + score_0_x527;
      res_1_sum <= res_1_sum + score_1_x527;
      res_2_sum <= res_2_sum + score_2_x527;
      res_3_sum <= res_3_sum + score_3_x527;
      res_4_sum <= res_4_sum + score_4_x527;
      res_5_sum <= res_5_sum + score_5_x527;
      res_6_sum <= res_6_sum + score_6_x527;
      res_7_sum <= res_7_sum + score_7_x527;
      res_8_sum <= res_8_sum + score_8_x527;
      res_9_sum <= res_9_sum + score_9_x527;
   end
   else if(res_done_x528) begin
      res_0_sum <= res_0_sum + score_0_x528;
      res_1_sum <= res_1_sum + score_1_x528;
      res_2_sum <= res_2_sum + score_2_x528;
      res_3_sum <= res_3_sum + score_3_x528;
      res_4_sum <= res_4_sum + score_4_x528;
      res_5_sum <= res_5_sum + score_5_x528;
      res_6_sum <= res_6_sum + score_6_x528;
      res_7_sum <= res_7_sum + score_7_x528;
      res_8_sum <= res_8_sum + score_8_x528;
      res_9_sum <= res_9_sum + score_9_x528;
   end
   else if(res_done_x529) begin
      res_0_sum <= res_0_sum + score_0_x529;
      res_1_sum <= res_1_sum + score_1_x529;
      res_2_sum <= res_2_sum + score_2_x529;
      res_3_sum <= res_3_sum + score_3_x529;
      res_4_sum <= res_4_sum + score_4_x529;
      res_5_sum <= res_5_sum + score_5_x529;
      res_6_sum <= res_6_sum + score_6_x529;
      res_7_sum <= res_7_sum + score_7_x529;
      res_8_sum <= res_8_sum + score_8_x529;
      res_9_sum <= res_9_sum + score_9_x529;
   end
   else if(res_done_x530) begin
      res_0_sum <= res_0_sum + score_0_x530;
      res_1_sum <= res_1_sum + score_1_x530;
      res_2_sum <= res_2_sum + score_2_x530;
      res_3_sum <= res_3_sum + score_3_x530;
      res_4_sum <= res_4_sum + score_4_x530;
      res_5_sum <= res_5_sum + score_5_x530;
      res_6_sum <= res_6_sum + score_6_x530;
      res_7_sum <= res_7_sum + score_7_x530;
      res_8_sum <= res_8_sum + score_8_x530;
      res_9_sum <= res_9_sum + score_9_x530;
   end
   else if(res_done_x531) begin
      res_0_sum <= res_0_sum + score_0_x531;
      res_1_sum <= res_1_sum + score_1_x531;
      res_2_sum <= res_2_sum + score_2_x531;
      res_3_sum <= res_3_sum + score_3_x531;
      res_4_sum <= res_4_sum + score_4_x531;
      res_5_sum <= res_5_sum + score_5_x531;
      res_6_sum <= res_6_sum + score_6_x531;
      res_7_sum <= res_7_sum + score_7_x531;
      res_8_sum <= res_8_sum + score_8_x531;
      res_9_sum <= res_9_sum + score_9_x531;
   end
   else if(res_done_x532) begin
      res_0_sum <= res_0_sum + score_0_x532;
      res_1_sum <= res_1_sum + score_1_x532;
      res_2_sum <= res_2_sum + score_2_x532;
      res_3_sum <= res_3_sum + score_3_x532;
      res_4_sum <= res_4_sum + score_4_x532;
      res_5_sum <= res_5_sum + score_5_x532;
      res_6_sum <= res_6_sum + score_6_x532;
      res_7_sum <= res_7_sum + score_7_x532;
      res_8_sum <= res_8_sum + score_8_x532;
      res_9_sum <= res_9_sum + score_9_x532;
   end
   else if(res_done_x533) begin
      res_0_sum <= res_0_sum + score_0_x533;
      res_1_sum <= res_1_sum + score_1_x533;
      res_2_sum <= res_2_sum + score_2_x533;
      res_3_sum <= res_3_sum + score_3_x533;
      res_4_sum <= res_4_sum + score_4_x533;
      res_5_sum <= res_5_sum + score_5_x533;
      res_6_sum <= res_6_sum + score_6_x533;
      res_7_sum <= res_7_sum + score_7_x533;
      res_8_sum <= res_8_sum + score_8_x533;
      res_9_sum <= res_9_sum + score_9_x533;
   end
   else if(res_done_x534) begin
      res_0_sum <= res_0_sum + score_0_x534;
      res_1_sum <= res_1_sum + score_1_x534;
      res_2_sum <= res_2_sum + score_2_x534;
      res_3_sum <= res_3_sum + score_3_x534;
      res_4_sum <= res_4_sum + score_4_x534;
      res_5_sum <= res_5_sum + score_5_x534;
      res_6_sum <= res_6_sum + score_6_x534;
      res_7_sum <= res_7_sum + score_7_x534;
      res_8_sum <= res_8_sum + score_8_x534;
      res_9_sum <= res_9_sum + score_9_x534;
   end
   else if(res_done_x535) begin
      res_0_sum <= res_0_sum + score_0_x535;
      res_1_sum <= res_1_sum + score_1_x535;
      res_2_sum <= res_2_sum + score_2_x535;
      res_3_sum <= res_3_sum + score_3_x535;
      res_4_sum <= res_4_sum + score_4_x535;
      res_5_sum <= res_5_sum + score_5_x535;
      res_6_sum <= res_6_sum + score_6_x535;
      res_7_sum <= res_7_sum + score_7_x535;
      res_8_sum <= res_8_sum + score_8_x535;
      res_9_sum <= res_9_sum + score_9_x535;
   end
   else if(res_done_x536) begin
      res_0_sum <= res_0_sum + score_0_x536;
      res_1_sum <= res_1_sum + score_1_x536;
      res_2_sum <= res_2_sum + score_2_x536;
      res_3_sum <= res_3_sum + score_3_x536;
      res_4_sum <= res_4_sum + score_4_x536;
      res_5_sum <= res_5_sum + score_5_x536;
      res_6_sum <= res_6_sum + score_6_x536;
      res_7_sum <= res_7_sum + score_7_x536;
      res_8_sum <= res_8_sum + score_8_x536;
      res_9_sum <= res_9_sum + score_9_x536;
   end
   else if(res_done_x537) begin
      res_0_sum <= res_0_sum + score_0_x537;
      res_1_sum <= res_1_sum + score_1_x537;
      res_2_sum <= res_2_sum + score_2_x537;
      res_3_sum <= res_3_sum + score_3_x537;
      res_4_sum <= res_4_sum + score_4_x537;
      res_5_sum <= res_5_sum + score_5_x537;
      res_6_sum <= res_6_sum + score_6_x537;
      res_7_sum <= res_7_sum + score_7_x537;
      res_8_sum <= res_8_sum + score_8_x537;
      res_9_sum <= res_9_sum + score_9_x537;
   end
   else if(res_done_x538) begin
      res_0_sum <= res_0_sum + score_0_x538;
      res_1_sum <= res_1_sum + score_1_x538;
      res_2_sum <= res_2_sum + score_2_x538;
      res_3_sum <= res_3_sum + score_3_x538;
      res_4_sum <= res_4_sum + score_4_x538;
      res_5_sum <= res_5_sum + score_5_x538;
      res_6_sum <= res_6_sum + score_6_x538;
      res_7_sum <= res_7_sum + score_7_x538;
      res_8_sum <= res_8_sum + score_8_x538;
      res_9_sum <= res_9_sum + score_9_x538;
   end
   else if(res_done_x539) begin
      res_0_sum <= res_0_sum + score_0_x539;
      res_1_sum <= res_1_sum + score_1_x539;
      res_2_sum <= res_2_sum + score_2_x539;
      res_3_sum <= res_3_sum + score_3_x539;
      res_4_sum <= res_4_sum + score_4_x539;
      res_5_sum <= res_5_sum + score_5_x539;
      res_6_sum <= res_6_sum + score_6_x539;
      res_7_sum <= res_7_sum + score_7_x539;
      res_8_sum <= res_8_sum + score_8_x539;
      res_9_sum <= res_9_sum + score_9_x539;
   end
   else if(res_done_x540) begin
      res_0_sum <= res_0_sum + score_0_x540;
      res_1_sum <= res_1_sum + score_1_x540;
      res_2_sum <= res_2_sum + score_2_x540;
      res_3_sum <= res_3_sum + score_3_x540;
      res_4_sum <= res_4_sum + score_4_x540;
      res_5_sum <= res_5_sum + score_5_x540;
      res_6_sum <= res_6_sum + score_6_x540;
      res_7_sum <= res_7_sum + score_7_x540;
      res_8_sum <= res_8_sum + score_8_x540;
      res_9_sum <= res_9_sum + score_9_x540;
   end
   else if(res_done_x541) begin
      res_0_sum <= res_0_sum + score_0_x541;
      res_1_sum <= res_1_sum + score_1_x541;
      res_2_sum <= res_2_sum + score_2_x541;
      res_3_sum <= res_3_sum + score_3_x541;
      res_4_sum <= res_4_sum + score_4_x541;
      res_5_sum <= res_5_sum + score_5_x541;
      res_6_sum <= res_6_sum + score_6_x541;
      res_7_sum <= res_7_sum + score_7_x541;
      res_8_sum <= res_8_sum + score_8_x541;
      res_9_sum <= res_9_sum + score_9_x541;
   end
   else if(res_done_x542) begin
      res_0_sum <= res_0_sum + score_0_x542;
      res_1_sum <= res_1_sum + score_1_x542;
      res_2_sum <= res_2_sum + score_2_x542;
      res_3_sum <= res_3_sum + score_3_x542;
      res_4_sum <= res_4_sum + score_4_x542;
      res_5_sum <= res_5_sum + score_5_x542;
      res_6_sum <= res_6_sum + score_6_x542;
      res_7_sum <= res_7_sum + score_7_x542;
      res_8_sum <= res_8_sum + score_8_x542;
      res_9_sum <= res_9_sum + score_9_x542;
   end
   else if(res_done_x543) begin
      res_0_sum <= res_0_sum + score_0_x543;
      res_1_sum <= res_1_sum + score_1_x543;
      res_2_sum <= res_2_sum + score_2_x543;
      res_3_sum <= res_3_sum + score_3_x543;
      res_4_sum <= res_4_sum + score_4_x543;
      res_5_sum <= res_5_sum + score_5_x543;
      res_6_sum <= res_6_sum + score_6_x543;
      res_7_sum <= res_7_sum + score_7_x543;
      res_8_sum <= res_8_sum + score_8_x543;
      res_9_sum <= res_9_sum + score_9_x543;
   end
   else if(res_done_x544) begin
      res_0_sum <= res_0_sum + score_0_x544;
      res_1_sum <= res_1_sum + score_1_x544;
      res_2_sum <= res_2_sum + score_2_x544;
      res_3_sum <= res_3_sum + score_3_x544;
      res_4_sum <= res_4_sum + score_4_x544;
      res_5_sum <= res_5_sum + score_5_x544;
      res_6_sum <= res_6_sum + score_6_x544;
      res_7_sum <= res_7_sum + score_7_x544;
      res_8_sum <= res_8_sum + score_8_x544;
      res_9_sum <= res_9_sum + score_9_x544;
   end
   else if(res_done_x545) begin
      res_0_sum <= res_0_sum + score_0_x545;
      res_1_sum <= res_1_sum + score_1_x545;
      res_2_sum <= res_2_sum + score_2_x545;
      res_3_sum <= res_3_sum + score_3_x545;
      res_4_sum <= res_4_sum + score_4_x545;
      res_5_sum <= res_5_sum + score_5_x545;
      res_6_sum <= res_6_sum + score_6_x545;
      res_7_sum <= res_7_sum + score_7_x545;
      res_8_sum <= res_8_sum + score_8_x545;
      res_9_sum <= res_9_sum + score_9_x545;
   end
   else if(res_done_x546) begin
      res_0_sum <= res_0_sum + score_0_x546;
      res_1_sum <= res_1_sum + score_1_x546;
      res_2_sum <= res_2_sum + score_2_x546;
      res_3_sum <= res_3_sum + score_3_x546;
      res_4_sum <= res_4_sum + score_4_x546;
      res_5_sum <= res_5_sum + score_5_x546;
      res_6_sum <= res_6_sum + score_6_x546;
      res_7_sum <= res_7_sum + score_7_x546;
      res_8_sum <= res_8_sum + score_8_x546;
      res_9_sum <= res_9_sum + score_9_x546;
   end
   else if(res_done_x547) begin
      res_0_sum <= res_0_sum + score_0_x547;
      res_1_sum <= res_1_sum + score_1_x547;
      res_2_sum <= res_2_sum + score_2_x547;
      res_3_sum <= res_3_sum + score_3_x547;
      res_4_sum <= res_4_sum + score_4_x547;
      res_5_sum <= res_5_sum + score_5_x547;
      res_6_sum <= res_6_sum + score_6_x547;
      res_7_sum <= res_7_sum + score_7_x547;
      res_8_sum <= res_8_sum + score_8_x547;
      res_9_sum <= res_9_sum + score_9_x547;
   end
   else if(res_done_x548) begin
      res_0_sum <= res_0_sum + score_0_x548;
      res_1_sum <= res_1_sum + score_1_x548;
      res_2_sum <= res_2_sum + score_2_x548;
      res_3_sum <= res_3_sum + score_3_x548;
      res_4_sum <= res_4_sum + score_4_x548;
      res_5_sum <= res_5_sum + score_5_x548;
      res_6_sum <= res_6_sum + score_6_x548;
      res_7_sum <= res_7_sum + score_7_x548;
      res_8_sum <= res_8_sum + score_8_x548;
      res_9_sum <= res_9_sum + score_9_x548;
   end
   else if(res_done_x549) begin
      res_0_sum <= res_0_sum + score_0_x549;
      res_1_sum <= res_1_sum + score_1_x549;
      res_2_sum <= res_2_sum + score_2_x549;
      res_3_sum <= res_3_sum + score_3_x549;
      res_4_sum <= res_4_sum + score_4_x549;
      res_5_sum <= res_5_sum + score_5_x549;
      res_6_sum <= res_6_sum + score_6_x549;
      res_7_sum <= res_7_sum + score_7_x549;
      res_8_sum <= res_8_sum + score_8_x549;
      res_9_sum <= res_9_sum + score_9_x549;
   end
   else if(res_done_x550) begin
      res_0_sum <= res_0_sum + score_0_x550;
      res_1_sum <= res_1_sum + score_1_x550;
      res_2_sum <= res_2_sum + score_2_x550;
      res_3_sum <= res_3_sum + score_3_x550;
      res_4_sum <= res_4_sum + score_4_x550;
      res_5_sum <= res_5_sum + score_5_x550;
      res_6_sum <= res_6_sum + score_6_x550;
      res_7_sum <= res_7_sum + score_7_x550;
      res_8_sum <= res_8_sum + score_8_x550;
      res_9_sum <= res_9_sum + score_9_x550;
   end
   else if(res_done_x551) begin
      res_0_sum <= res_0_sum + score_0_x551;
      res_1_sum <= res_1_sum + score_1_x551;
      res_2_sum <= res_2_sum + score_2_x551;
      res_3_sum <= res_3_sum + score_3_x551;
      res_4_sum <= res_4_sum + score_4_x551;
      res_5_sum <= res_5_sum + score_5_x551;
      res_6_sum <= res_6_sum + score_6_x551;
      res_7_sum <= res_7_sum + score_7_x551;
      res_8_sum <= res_8_sum + score_8_x551;
      res_9_sum <= res_9_sum + score_9_x551;
   end
   else if(res_done_x552) begin
      res_0_sum <= res_0_sum + score_0_x552;
      res_1_sum <= res_1_sum + score_1_x552;
      res_2_sum <= res_2_sum + score_2_x552;
      res_3_sum <= res_3_sum + score_3_x552;
      res_4_sum <= res_4_sum + score_4_x552;
      res_5_sum <= res_5_sum + score_5_x552;
      res_6_sum <= res_6_sum + score_6_x552;
      res_7_sum <= res_7_sum + score_7_x552;
      res_8_sum <= res_8_sum + score_8_x552;
      res_9_sum <= res_9_sum + score_9_x552;
   end
   else if(res_done_x553) begin
      res_0_sum <= res_0_sum + score_0_x553;
      res_1_sum <= res_1_sum + score_1_x553;
      res_2_sum <= res_2_sum + score_2_x553;
      res_3_sum <= res_3_sum + score_3_x553;
      res_4_sum <= res_4_sum + score_4_x553;
      res_5_sum <= res_5_sum + score_5_x553;
      res_6_sum <= res_6_sum + score_6_x553;
      res_7_sum <= res_7_sum + score_7_x553;
      res_8_sum <= res_8_sum + score_8_x553;
      res_9_sum <= res_9_sum + score_9_x553;
   end
   else if(res_done_x554) begin
      res_0_sum <= res_0_sum + score_0_x554;
      res_1_sum <= res_1_sum + score_1_x554;
      res_2_sum <= res_2_sum + score_2_x554;
      res_3_sum <= res_3_sum + score_3_x554;
      res_4_sum <= res_4_sum + score_4_x554;
      res_5_sum <= res_5_sum + score_5_x554;
      res_6_sum <= res_6_sum + score_6_x554;
      res_7_sum <= res_7_sum + score_7_x554;
      res_8_sum <= res_8_sum + score_8_x554;
      res_9_sum <= res_9_sum + score_9_x554;
   end
   else if(res_done_x555) begin
      res_0_sum <= res_0_sum + score_0_x555;
      res_1_sum <= res_1_sum + score_1_x555;
      res_2_sum <= res_2_sum + score_2_x555;
      res_3_sum <= res_3_sum + score_3_x555;
      res_4_sum <= res_4_sum + score_4_x555;
      res_5_sum <= res_5_sum + score_5_x555;
      res_6_sum <= res_6_sum + score_6_x555;
      res_7_sum <= res_7_sum + score_7_x555;
      res_8_sum <= res_8_sum + score_8_x555;
      res_9_sum <= res_9_sum + score_9_x555;
   end
   else if(res_done_x556) begin
      res_0_sum <= res_0_sum + score_0_x556;
      res_1_sum <= res_1_sum + score_1_x556;
      res_2_sum <= res_2_sum + score_2_x556;
      res_3_sum <= res_3_sum + score_3_x556;
      res_4_sum <= res_4_sum + score_4_x556;
      res_5_sum <= res_5_sum + score_5_x556;
      res_6_sum <= res_6_sum + score_6_x556;
      res_7_sum <= res_7_sum + score_7_x556;
      res_8_sum <= res_8_sum + score_8_x556;
      res_9_sum <= res_9_sum + score_9_x556;
   end
   else if(res_done_x557) begin
      res_0_sum <= res_0_sum + score_0_x557;
      res_1_sum <= res_1_sum + score_1_x557;
      res_2_sum <= res_2_sum + score_2_x557;
      res_3_sum <= res_3_sum + score_3_x557;
      res_4_sum <= res_4_sum + score_4_x557;
      res_5_sum <= res_5_sum + score_5_x557;
      res_6_sum <= res_6_sum + score_6_x557;
      res_7_sum <= res_7_sum + score_7_x557;
      res_8_sum <= res_8_sum + score_8_x557;
      res_9_sum <= res_9_sum + score_9_x557;
   end
   else if(res_done_x558) begin
      res_0_sum <= res_0_sum + score_0_x558;
      res_1_sum <= res_1_sum + score_1_x558;
      res_2_sum <= res_2_sum + score_2_x558;
      res_3_sum <= res_3_sum + score_3_x558;
      res_4_sum <= res_4_sum + score_4_x558;
      res_5_sum <= res_5_sum + score_5_x558;
      res_6_sum <= res_6_sum + score_6_x558;
      res_7_sum <= res_7_sum + score_7_x558;
      res_8_sum <= res_8_sum + score_8_x558;
      res_9_sum <= res_9_sum + score_9_x558;
   end
   else if(res_done_x559) begin
      res_0_sum <= res_0_sum + score_0_x559;
      res_1_sum <= res_1_sum + score_1_x559;
      res_2_sum <= res_2_sum + score_2_x559;
      res_3_sum <= res_3_sum + score_3_x559;
      res_4_sum <= res_4_sum + score_4_x559;
      res_5_sum <= res_5_sum + score_5_x559;
      res_6_sum <= res_6_sum + score_6_x559;
      res_7_sum <= res_7_sum + score_7_x559;
      res_8_sum <= res_8_sum + score_8_x559;
      res_9_sum <= res_9_sum + score_9_x559;
   end
   else if(res_done_x560) begin
      res_0_sum <= res_0_sum + score_0_x560;
      res_1_sum <= res_1_sum + score_1_x560;
      res_2_sum <= res_2_sum + score_2_x560;
      res_3_sum <= res_3_sum + score_3_x560;
      res_4_sum <= res_4_sum + score_4_x560;
      res_5_sum <= res_5_sum + score_5_x560;
      res_6_sum <= res_6_sum + score_6_x560;
      res_7_sum <= res_7_sum + score_7_x560;
      res_8_sum <= res_8_sum + score_8_x560;
      res_9_sum <= res_9_sum + score_9_x560;
   end
   else if(res_done_x561) begin
      res_0_sum <= res_0_sum + score_0_x561;
      res_1_sum <= res_1_sum + score_1_x561;
      res_2_sum <= res_2_sum + score_2_x561;
      res_3_sum <= res_3_sum + score_3_x561;
      res_4_sum <= res_4_sum + score_4_x561;
      res_5_sum <= res_5_sum + score_5_x561;
      res_6_sum <= res_6_sum + score_6_x561;
      res_7_sum <= res_7_sum + score_7_x561;
      res_8_sum <= res_8_sum + score_8_x561;
      res_9_sum <= res_9_sum + score_9_x561;
   end
   else if(res_done_x562) begin
      res_0_sum <= res_0_sum + score_0_x562;
      res_1_sum <= res_1_sum + score_1_x562;
      res_2_sum <= res_2_sum + score_2_x562;
      res_3_sum <= res_3_sum + score_3_x562;
      res_4_sum <= res_4_sum + score_4_x562;
      res_5_sum <= res_5_sum + score_5_x562;
      res_6_sum <= res_6_sum + score_6_x562;
      res_7_sum <= res_7_sum + score_7_x562;
      res_8_sum <= res_8_sum + score_8_x562;
      res_9_sum <= res_9_sum + score_9_x562;
   end
   else if(res_done_x563) begin
      res_0_sum <= res_0_sum + score_0_x563;
      res_1_sum <= res_1_sum + score_1_x563;
      res_2_sum <= res_2_sum + score_2_x563;
      res_3_sum <= res_3_sum + score_3_x563;
      res_4_sum <= res_4_sum + score_4_x563;
      res_5_sum <= res_5_sum + score_5_x563;
      res_6_sum <= res_6_sum + score_6_x563;
      res_7_sum <= res_7_sum + score_7_x563;
      res_8_sum <= res_8_sum + score_8_x563;
      res_9_sum <= res_9_sum + score_9_x563;
   end
   else if(res_done_x564) begin
      res_0_sum <= res_0_sum + score_0_x564;
      res_1_sum <= res_1_sum + score_1_x564;
      res_2_sum <= res_2_sum + score_2_x564;
      res_3_sum <= res_3_sum + score_3_x564;
      res_4_sum <= res_4_sum + score_4_x564;
      res_5_sum <= res_5_sum + score_5_x564;
      res_6_sum <= res_6_sum + score_6_x564;
      res_7_sum <= res_7_sum + score_7_x564;
      res_8_sum <= res_8_sum + score_8_x564;
      res_9_sum <= res_9_sum + score_9_x564;
   end
   else if(res_done_x565) begin
      res_0_sum <= res_0_sum + score_0_x565;
      res_1_sum <= res_1_sum + score_1_x565;
      res_2_sum <= res_2_sum + score_2_x565;
      res_3_sum <= res_3_sum + score_3_x565;
      res_4_sum <= res_4_sum + score_4_x565;
      res_5_sum <= res_5_sum + score_5_x565;
      res_6_sum <= res_6_sum + score_6_x565;
      res_7_sum <= res_7_sum + score_7_x565;
      res_8_sum <= res_8_sum + score_8_x565;
      res_9_sum <= res_9_sum + score_9_x565;
   end
   else if(res_done_x566) begin
      res_0_sum <= res_0_sum + score_0_x566;
      res_1_sum <= res_1_sum + score_1_x566;
      res_2_sum <= res_2_sum + score_2_x566;
      res_3_sum <= res_3_sum + score_3_x566;
      res_4_sum <= res_4_sum + score_4_x566;
      res_5_sum <= res_5_sum + score_5_x566;
      res_6_sum <= res_6_sum + score_6_x566;
      res_7_sum <= res_7_sum + score_7_x566;
      res_8_sum <= res_8_sum + score_8_x566;
      res_9_sum <= res_9_sum + score_9_x566;
   end
   else if(res_done_x567) begin
      res_0_sum <= res_0_sum + score_0_x567;
      res_1_sum <= res_1_sum + score_1_x567;
      res_2_sum <= res_2_sum + score_2_x567;
      res_3_sum <= res_3_sum + score_3_x567;
      res_4_sum <= res_4_sum + score_4_x567;
      res_5_sum <= res_5_sum + score_5_x567;
      res_6_sum <= res_6_sum + score_6_x567;
      res_7_sum <= res_7_sum + score_7_x567;
      res_8_sum <= res_8_sum + score_8_x567;
      res_9_sum <= res_9_sum + score_9_x567;
   end
   else if(res_done_x568) begin
      res_0_sum <= res_0_sum + score_0_x568;
      res_1_sum <= res_1_sum + score_1_x568;
      res_2_sum <= res_2_sum + score_2_x568;
      res_3_sum <= res_3_sum + score_3_x568;
      res_4_sum <= res_4_sum + score_4_x568;
      res_5_sum <= res_5_sum + score_5_x568;
      res_6_sum <= res_6_sum + score_6_x568;
      res_7_sum <= res_7_sum + score_7_x568;
      res_8_sum <= res_8_sum + score_8_x568;
      res_9_sum <= res_9_sum + score_9_x568;
   end
   else if(res_done_x569) begin
      res_0_sum <= res_0_sum + score_0_x569;
      res_1_sum <= res_1_sum + score_1_x569;
      res_2_sum <= res_2_sum + score_2_x569;
      res_3_sum <= res_3_sum + score_3_x569;
      res_4_sum <= res_4_sum + score_4_x569;
      res_5_sum <= res_5_sum + score_5_x569;
      res_6_sum <= res_6_sum + score_6_x569;
      res_7_sum <= res_7_sum + score_7_x569;
      res_8_sum <= res_8_sum + score_8_x569;
      res_9_sum <= res_9_sum + score_9_x569;
   end
   else if(res_done_x570) begin
      res_0_sum <= res_0_sum + score_0_x570;
      res_1_sum <= res_1_sum + score_1_x570;
      res_2_sum <= res_2_sum + score_2_x570;
      res_3_sum <= res_3_sum + score_3_x570;
      res_4_sum <= res_4_sum + score_4_x570;
      res_5_sum <= res_5_sum + score_5_x570;
      res_6_sum <= res_6_sum + score_6_x570;
      res_7_sum <= res_7_sum + score_7_x570;
      res_8_sum <= res_8_sum + score_8_x570;
      res_9_sum <= res_9_sum + score_9_x570;
   end
   else if(res_done_x571) begin
      res_0_sum <= res_0_sum + score_0_x571;
      res_1_sum <= res_1_sum + score_1_x571;
      res_2_sum <= res_2_sum + score_2_x571;
      res_3_sum <= res_3_sum + score_3_x571;
      res_4_sum <= res_4_sum + score_4_x571;
      res_5_sum <= res_5_sum + score_5_x571;
      res_6_sum <= res_6_sum + score_6_x571;
      res_7_sum <= res_7_sum + score_7_x571;
      res_8_sum <= res_8_sum + score_8_x571;
      res_9_sum <= res_9_sum + score_9_x571;
   end
   else if(res_done_x572) begin
      res_0_sum <= res_0_sum + score_0_x572;
      res_1_sum <= res_1_sum + score_1_x572;
      res_2_sum <= res_2_sum + score_2_x572;
      res_3_sum <= res_3_sum + score_3_x572;
      res_4_sum <= res_4_sum + score_4_x572;
      res_5_sum <= res_5_sum + score_5_x572;
      res_6_sum <= res_6_sum + score_6_x572;
      res_7_sum <= res_7_sum + score_7_x572;
      res_8_sum <= res_8_sum + score_8_x572;
      res_9_sum <= res_9_sum + score_9_x572;
   end
   else if(res_done_x573) begin
      res_0_sum <= res_0_sum + score_0_x573;
      res_1_sum <= res_1_sum + score_1_x573;
      res_2_sum <= res_2_sum + score_2_x573;
      res_3_sum <= res_3_sum + score_3_x573;
      res_4_sum <= res_4_sum + score_4_x573;
      res_5_sum <= res_5_sum + score_5_x573;
      res_6_sum <= res_6_sum + score_6_x573;
      res_7_sum <= res_7_sum + score_7_x573;
      res_8_sum <= res_8_sum + score_8_x573;
      res_9_sum <= res_9_sum + score_9_x573;
   end
   else if(res_done_x574) begin
      res_0_sum <= res_0_sum + score_0_x574;
      res_1_sum <= res_1_sum + score_1_x574;
      res_2_sum <= res_2_sum + score_2_x574;
      res_3_sum <= res_3_sum + score_3_x574;
      res_4_sum <= res_4_sum + score_4_x574;
      res_5_sum <= res_5_sum + score_5_x574;
      res_6_sum <= res_6_sum + score_6_x574;
      res_7_sum <= res_7_sum + score_7_x574;
      res_8_sum <= res_8_sum + score_8_x574;
      res_9_sum <= res_9_sum + score_9_x574;
   end
   else if(res_done_x575) begin
      res_0_sum <= res_0_sum + score_0_x575;
      res_1_sum <= res_1_sum + score_1_x575;
      res_2_sum <= res_2_sum + score_2_x575;
      res_3_sum <= res_3_sum + score_3_x575;
      res_4_sum <= res_4_sum + score_4_x575;
      res_5_sum <= res_5_sum + score_5_x575;
      res_6_sum <= res_6_sum + score_6_x575;
      res_7_sum <= res_7_sum + score_7_x575;
      res_8_sum <= res_8_sum + score_8_x575;
      res_9_sum <= res_9_sum + score_9_x575;
   end
   else if(res_done_x576) begin
      res_0_sum <= res_0_sum + score_0_x576;
      res_1_sum <= res_1_sum + score_1_x576;
      res_2_sum <= res_2_sum + score_2_x576;
      res_3_sum <= res_3_sum + score_3_x576;
      res_4_sum <= res_4_sum + score_4_x576;
      res_5_sum <= res_5_sum + score_5_x576;
      res_6_sum <= res_6_sum + score_6_x576;
      res_7_sum <= res_7_sum + score_7_x576;
      res_8_sum <= res_8_sum + score_8_x576;
      res_9_sum <= res_9_sum + score_9_x576;
   end
   else if(res_done_x577) begin
      res_0_sum <= res_0_sum + score_0_x577;
      res_1_sum <= res_1_sum + score_1_x577;
      res_2_sum <= res_2_sum + score_2_x577;
      res_3_sum <= res_3_sum + score_3_x577;
      res_4_sum <= res_4_sum + score_4_x577;
      res_5_sum <= res_5_sum + score_5_x577;
      res_6_sum <= res_6_sum + score_6_x577;
      res_7_sum <= res_7_sum + score_7_x577;
      res_8_sum <= res_8_sum + score_8_x577;
      res_9_sum <= res_9_sum + score_9_x577;
   end
   else if(res_done_x578) begin
      res_0_sum <= res_0_sum + score_0_x578;
      res_1_sum <= res_1_sum + score_1_x578;
      res_2_sum <= res_2_sum + score_2_x578;
      res_3_sum <= res_3_sum + score_3_x578;
      res_4_sum <= res_4_sum + score_4_x578;
      res_5_sum <= res_5_sum + score_5_x578;
      res_6_sum <= res_6_sum + score_6_x578;
      res_7_sum <= res_7_sum + score_7_x578;
      res_8_sum <= res_8_sum + score_8_x578;
      res_9_sum <= res_9_sum + score_9_x578;
   end
   else if(res_done_x579) begin
      res_0_sum <= res_0_sum + score_0_x579;
      res_1_sum <= res_1_sum + score_1_x579;
      res_2_sum <= res_2_sum + score_2_x579;
      res_3_sum <= res_3_sum + score_3_x579;
      res_4_sum <= res_4_sum + score_4_x579;
      res_5_sum <= res_5_sum + score_5_x579;
      res_6_sum <= res_6_sum + score_6_x579;
      res_7_sum <= res_7_sum + score_7_x579;
      res_8_sum <= res_8_sum + score_8_x579;
      res_9_sum <= res_9_sum + score_9_x579;
   end
   else if(res_done_x580) begin
      res_0_sum <= res_0_sum + score_0_x580;
      res_1_sum <= res_1_sum + score_1_x580;
      res_2_sum <= res_2_sum + score_2_x580;
      res_3_sum <= res_3_sum + score_3_x580;
      res_4_sum <= res_4_sum + score_4_x580;
      res_5_sum <= res_5_sum + score_5_x580;
      res_6_sum <= res_6_sum + score_6_x580;
      res_7_sum <= res_7_sum + score_7_x580;
      res_8_sum <= res_8_sum + score_8_x580;
      res_9_sum <= res_9_sum + score_9_x580;
   end
   else if(res_done_x581) begin
      res_0_sum <= res_0_sum + score_0_x581;
      res_1_sum <= res_1_sum + score_1_x581;
      res_2_sum <= res_2_sum + score_2_x581;
      res_3_sum <= res_3_sum + score_3_x581;
      res_4_sum <= res_4_sum + score_4_x581;
      res_5_sum <= res_5_sum + score_5_x581;
      res_6_sum <= res_6_sum + score_6_x581;
      res_7_sum <= res_7_sum + score_7_x581;
      res_8_sum <= res_8_sum + score_8_x581;
      res_9_sum <= res_9_sum + score_9_x581;
   end
   else if(res_done_x582) begin
      res_0_sum <= res_0_sum + score_0_x582;
      res_1_sum <= res_1_sum + score_1_x582;
      res_2_sum <= res_2_sum + score_2_x582;
      res_3_sum <= res_3_sum + score_3_x582;
      res_4_sum <= res_4_sum + score_4_x582;
      res_5_sum <= res_5_sum + score_5_x582;
      res_6_sum <= res_6_sum + score_6_x582;
      res_7_sum <= res_7_sum + score_7_x582;
      res_8_sum <= res_8_sum + score_8_x582;
      res_9_sum <= res_9_sum + score_9_x582;
   end
   else if(res_done_x583) begin
      res_0_sum <= res_0_sum + score_0_x583;
      res_1_sum <= res_1_sum + score_1_x583;
      res_2_sum <= res_2_sum + score_2_x583;
      res_3_sum <= res_3_sum + score_3_x583;
      res_4_sum <= res_4_sum + score_4_x583;
      res_5_sum <= res_5_sum + score_5_x583;
      res_6_sum <= res_6_sum + score_6_x583;
      res_7_sum <= res_7_sum + score_7_x583;
      res_8_sum <= res_8_sum + score_8_x583;
      res_9_sum <= res_9_sum + score_9_x583;
   end
   else if(res_done_x584) begin
      res_0_sum <= res_0_sum + score_0_x584;
      res_1_sum <= res_1_sum + score_1_x584;
      res_2_sum <= res_2_sum + score_2_x584;
      res_3_sum <= res_3_sum + score_3_x584;
      res_4_sum <= res_4_sum + score_4_x584;
      res_5_sum <= res_5_sum + score_5_x584;
      res_6_sum <= res_6_sum + score_6_x584;
      res_7_sum <= res_7_sum + score_7_x584;
      res_8_sum <= res_8_sum + score_8_x584;
      res_9_sum <= res_9_sum + score_9_x584;
   end
   else if(res_done_x585) begin
      res_0_sum <= res_0_sum + score_0_x585;
      res_1_sum <= res_1_sum + score_1_x585;
      res_2_sum <= res_2_sum + score_2_x585;
      res_3_sum <= res_3_sum + score_3_x585;
      res_4_sum <= res_4_sum + score_4_x585;
      res_5_sum <= res_5_sum + score_5_x585;
      res_6_sum <= res_6_sum + score_6_x585;
      res_7_sum <= res_7_sum + score_7_x585;
      res_8_sum <= res_8_sum + score_8_x585;
      res_9_sum <= res_9_sum + score_9_x585;
   end
   else if(res_done_x586) begin
      res_0_sum <= res_0_sum + score_0_x586;
      res_1_sum <= res_1_sum + score_1_x586;
      res_2_sum <= res_2_sum + score_2_x586;
      res_3_sum <= res_3_sum + score_3_x586;
      res_4_sum <= res_4_sum + score_4_x586;
      res_5_sum <= res_5_sum + score_5_x586;
      res_6_sum <= res_6_sum + score_6_x586;
      res_7_sum <= res_7_sum + score_7_x586;
      res_8_sum <= res_8_sum + score_8_x586;
      res_9_sum <= res_9_sum + score_9_x586;
   end
   else if(res_done_x587) begin
      res_0_sum <= res_0_sum + score_0_x587;
      res_1_sum <= res_1_sum + score_1_x587;
      res_2_sum <= res_2_sum + score_2_x587;
      res_3_sum <= res_3_sum + score_3_x587;
      res_4_sum <= res_4_sum + score_4_x587;
      res_5_sum <= res_5_sum + score_5_x587;
      res_6_sum <= res_6_sum + score_6_x587;
      res_7_sum <= res_7_sum + score_7_x587;
      res_8_sum <= res_8_sum + score_8_x587;
      res_9_sum <= res_9_sum + score_9_x587;
   end
   else if(res_done_x588) begin
      res_0_sum <= res_0_sum + score_0_x588;
      res_1_sum <= res_1_sum + score_1_x588;
      res_2_sum <= res_2_sum + score_2_x588;
      res_3_sum <= res_3_sum + score_3_x588;
      res_4_sum <= res_4_sum + score_4_x588;
      res_5_sum <= res_5_sum + score_5_x588;
      res_6_sum <= res_6_sum + score_6_x588;
      res_7_sum <= res_7_sum + score_7_x588;
      res_8_sum <= res_8_sum + score_8_x588;
      res_9_sum <= res_9_sum + score_9_x588;
   end
   else if(res_done_x589) begin
      res_0_sum <= res_0_sum + score_0_x589;
      res_1_sum <= res_1_sum + score_1_x589;
      res_2_sum <= res_2_sum + score_2_x589;
      res_3_sum <= res_3_sum + score_3_x589;
      res_4_sum <= res_4_sum + score_4_x589;
      res_5_sum <= res_5_sum + score_5_x589;
      res_6_sum <= res_6_sum + score_6_x589;
      res_7_sum <= res_7_sum + score_7_x589;
      res_8_sum <= res_8_sum + score_8_x589;
      res_9_sum <= res_9_sum + score_9_x589;
   end
   else if(res_done_x590) begin
      res_0_sum <= res_0_sum + score_0_x590;
      res_1_sum <= res_1_sum + score_1_x590;
      res_2_sum <= res_2_sum + score_2_x590;
      res_3_sum <= res_3_sum + score_3_x590;
      res_4_sum <= res_4_sum + score_4_x590;
      res_5_sum <= res_5_sum + score_5_x590;
      res_6_sum <= res_6_sum + score_6_x590;
      res_7_sum <= res_7_sum + score_7_x590;
      res_8_sum <= res_8_sum + score_8_x590;
      res_9_sum <= res_9_sum + score_9_x590;
   end
   else if(res_done_x591) begin
      res_0_sum <= res_0_sum + score_0_x591;
      res_1_sum <= res_1_sum + score_1_x591;
      res_2_sum <= res_2_sum + score_2_x591;
      res_3_sum <= res_3_sum + score_3_x591;
      res_4_sum <= res_4_sum + score_4_x591;
      res_5_sum <= res_5_sum + score_5_x591;
      res_6_sum <= res_6_sum + score_6_x591;
      res_7_sum <= res_7_sum + score_7_x591;
      res_8_sum <= res_8_sum + score_8_x591;
      res_9_sum <= res_9_sum + score_9_x591;
   end
   else if(res_done_x592) begin
      res_0_sum <= res_0_sum + score_0_x592;
      res_1_sum <= res_1_sum + score_1_x592;
      res_2_sum <= res_2_sum + score_2_x592;
      res_3_sum <= res_3_sum + score_3_x592;
      res_4_sum <= res_4_sum + score_4_x592;
      res_5_sum <= res_5_sum + score_5_x592;
      res_6_sum <= res_6_sum + score_6_x592;
      res_7_sum <= res_7_sum + score_7_x592;
      res_8_sum <= res_8_sum + score_8_x592;
      res_9_sum <= res_9_sum + score_9_x592;
   end
   else if(res_done_x593) begin
      res_0_sum <= res_0_sum + score_0_x593;
      res_1_sum <= res_1_sum + score_1_x593;
      res_2_sum <= res_2_sum + score_2_x593;
      res_3_sum <= res_3_sum + score_3_x593;
      res_4_sum <= res_4_sum + score_4_x593;
      res_5_sum <= res_5_sum + score_5_x593;
      res_6_sum <= res_6_sum + score_6_x593;
      res_7_sum <= res_7_sum + score_7_x593;
      res_8_sum <= res_8_sum + score_8_x593;
      res_9_sum <= res_9_sum + score_9_x593;
   end
   else if(res_done_x594) begin
      res_0_sum <= res_0_sum + score_0_x594;
      res_1_sum <= res_1_sum + score_1_x594;
      res_2_sum <= res_2_sum + score_2_x594;
      res_3_sum <= res_3_sum + score_3_x594;
      res_4_sum <= res_4_sum + score_4_x594;
      res_5_sum <= res_5_sum + score_5_x594;
      res_6_sum <= res_6_sum + score_6_x594;
      res_7_sum <= res_7_sum + score_7_x594;
      res_8_sum <= res_8_sum + score_8_x594;
      res_9_sum <= res_9_sum + score_9_x594;
   end
   else if(res_done_x595) begin
      res_0_sum <= res_0_sum + score_0_x595;
      res_1_sum <= res_1_sum + score_1_x595;
      res_2_sum <= res_2_sum + score_2_x595;
      res_3_sum <= res_3_sum + score_3_x595;
      res_4_sum <= res_4_sum + score_4_x595;
      res_5_sum <= res_5_sum + score_5_x595;
      res_6_sum <= res_6_sum + score_6_x595;
      res_7_sum <= res_7_sum + score_7_x595;
      res_8_sum <= res_8_sum + score_8_x595;
      res_9_sum <= res_9_sum + score_9_x595;
   end
   else if(res_done_x596) begin
      res_0_sum <= res_0_sum + score_0_x596;
      res_1_sum <= res_1_sum + score_1_x596;
      res_2_sum <= res_2_sum + score_2_x596;
      res_3_sum <= res_3_sum + score_3_x596;
      res_4_sum <= res_4_sum + score_4_x596;
      res_5_sum <= res_5_sum + score_5_x596;
      res_6_sum <= res_6_sum + score_6_x596;
      res_7_sum <= res_7_sum + score_7_x596;
      res_8_sum <= res_8_sum + score_8_x596;
      res_9_sum <= res_9_sum + score_9_x596;
   end
   else if(res_done_x597) begin
      res_0_sum <= res_0_sum + score_0_x597;
      res_1_sum <= res_1_sum + score_1_x597;
      res_2_sum <= res_2_sum + score_2_x597;
      res_3_sum <= res_3_sum + score_3_x597;
      res_4_sum <= res_4_sum + score_4_x597;
      res_5_sum <= res_5_sum + score_5_x597;
      res_6_sum <= res_6_sum + score_6_x597;
      res_7_sum <= res_7_sum + score_7_x597;
      res_8_sum <= res_8_sum + score_8_x597;
      res_9_sum <= res_9_sum + score_9_x597;
   end
   else if(res_done_x598) begin
      res_0_sum <= res_0_sum + score_0_x598;
      res_1_sum <= res_1_sum + score_1_x598;
      res_2_sum <= res_2_sum + score_2_x598;
      res_3_sum <= res_3_sum + score_3_x598;
      res_4_sum <= res_4_sum + score_4_x598;
      res_5_sum <= res_5_sum + score_5_x598;
      res_6_sum <= res_6_sum + score_6_x598;
      res_7_sum <= res_7_sum + score_7_x598;
      res_8_sum <= res_8_sum + score_8_x598;
      res_9_sum <= res_9_sum + score_9_x598;
   end
   else if(res_done_x599) begin
      res_0_sum <= res_0_sum + score_0_x599;
      res_1_sum <= res_1_sum + score_1_x599;
      res_2_sum <= res_2_sum + score_2_x599;
      res_3_sum <= res_3_sum + score_3_x599;
      res_4_sum <= res_4_sum + score_4_x599;
      res_5_sum <= res_5_sum + score_5_x599;
      res_6_sum <= res_6_sum + score_6_x599;
      res_7_sum <= res_7_sum + score_7_x599;
      res_8_sum <= res_8_sum + score_8_x599;
      res_9_sum <= res_9_sum + score_9_x599;
   end
   else if(res_done_x600) begin
      res_0_sum <= res_0_sum + score_0_x600;
      res_1_sum <= res_1_sum + score_1_x600;
      res_2_sum <= res_2_sum + score_2_x600;
      res_3_sum <= res_3_sum + score_3_x600;
      res_4_sum <= res_4_sum + score_4_x600;
      res_5_sum <= res_5_sum + score_5_x600;
      res_6_sum <= res_6_sum + score_6_x600;
      res_7_sum <= res_7_sum + score_7_x600;
      res_8_sum <= res_8_sum + score_8_x600;
      res_9_sum <= res_9_sum + score_9_x600;
   end
   else if(res_done_x601) begin
      res_0_sum <= res_0_sum + score_0_x601;
      res_1_sum <= res_1_sum + score_1_x601;
      res_2_sum <= res_2_sum + score_2_x601;
      res_3_sum <= res_3_sum + score_3_x601;
      res_4_sum <= res_4_sum + score_4_x601;
      res_5_sum <= res_5_sum + score_5_x601;
      res_6_sum <= res_6_sum + score_6_x601;
      res_7_sum <= res_7_sum + score_7_x601;
      res_8_sum <= res_8_sum + score_8_x601;
      res_9_sum <= res_9_sum + score_9_x601;
   end
   else if(res_done_x602) begin
      res_0_sum <= res_0_sum + score_0_x602;
      res_1_sum <= res_1_sum + score_1_x602;
      res_2_sum <= res_2_sum + score_2_x602;
      res_3_sum <= res_3_sum + score_3_x602;
      res_4_sum <= res_4_sum + score_4_x602;
      res_5_sum <= res_5_sum + score_5_x602;
      res_6_sum <= res_6_sum + score_6_x602;
      res_7_sum <= res_7_sum + score_7_x602;
      res_8_sum <= res_8_sum + score_8_x602;
      res_9_sum <= res_9_sum + score_9_x602;
   end
   else if(res_done_x603) begin
      res_0_sum <= res_0_sum + score_0_x603;
      res_1_sum <= res_1_sum + score_1_x603;
      res_2_sum <= res_2_sum + score_2_x603;
      res_3_sum <= res_3_sum + score_3_x603;
      res_4_sum <= res_4_sum + score_4_x603;
      res_5_sum <= res_5_sum + score_5_x603;
      res_6_sum <= res_6_sum + score_6_x603;
      res_7_sum <= res_7_sum + score_7_x603;
      res_8_sum <= res_8_sum + score_8_x603;
      res_9_sum <= res_9_sum + score_9_x603;
   end
   else if(res_done_x604) begin
      res_0_sum <= res_0_sum + score_0_x604;
      res_1_sum <= res_1_sum + score_1_x604;
      res_2_sum <= res_2_sum + score_2_x604;
      res_3_sum <= res_3_sum + score_3_x604;
      res_4_sum <= res_4_sum + score_4_x604;
      res_5_sum <= res_5_sum + score_5_x604;
      res_6_sum <= res_6_sum + score_6_x604;
      res_7_sum <= res_7_sum + score_7_x604;
      res_8_sum <= res_8_sum + score_8_x604;
      res_9_sum <= res_9_sum + score_9_x604;
   end
   else if(res_done_x605) begin
      res_0_sum <= res_0_sum + score_0_x605;
      res_1_sum <= res_1_sum + score_1_x605;
      res_2_sum <= res_2_sum + score_2_x605;
      res_3_sum <= res_3_sum + score_3_x605;
      res_4_sum <= res_4_sum + score_4_x605;
      res_5_sum <= res_5_sum + score_5_x605;
      res_6_sum <= res_6_sum + score_6_x605;
      res_7_sum <= res_7_sum + score_7_x605;
      res_8_sum <= res_8_sum + score_8_x605;
      res_9_sum <= res_9_sum + score_9_x605;
   end
   else if(res_done_x606) begin
      res_0_sum <= res_0_sum + score_0_x606;
      res_1_sum <= res_1_sum + score_1_x606;
      res_2_sum <= res_2_sum + score_2_x606;
      res_3_sum <= res_3_sum + score_3_x606;
      res_4_sum <= res_4_sum + score_4_x606;
      res_5_sum <= res_5_sum + score_5_x606;
      res_6_sum <= res_6_sum + score_6_x606;
      res_7_sum <= res_7_sum + score_7_x606;
      res_8_sum <= res_8_sum + score_8_x606;
      res_9_sum <= res_9_sum + score_9_x606;
   end
   else if(res_done_x607) begin
      res_0_sum <= res_0_sum + score_0_x607;
      res_1_sum <= res_1_sum + score_1_x607;
      res_2_sum <= res_2_sum + score_2_x607;
      res_3_sum <= res_3_sum + score_3_x607;
      res_4_sum <= res_4_sum + score_4_x607;
      res_5_sum <= res_5_sum + score_5_x607;
      res_6_sum <= res_6_sum + score_6_x607;
      res_7_sum <= res_7_sum + score_7_x607;
      res_8_sum <= res_8_sum + score_8_x607;
      res_9_sum <= res_9_sum + score_9_x607;
   end
   else if(res_done_x608) begin
      res_0_sum <= res_0_sum + score_0_x608;
      res_1_sum <= res_1_sum + score_1_x608;
      res_2_sum <= res_2_sum + score_2_x608;
      res_3_sum <= res_3_sum + score_3_x608;
      res_4_sum <= res_4_sum + score_4_x608;
      res_5_sum <= res_5_sum + score_5_x608;
      res_6_sum <= res_6_sum + score_6_x608;
      res_7_sum <= res_7_sum + score_7_x608;
      res_8_sum <= res_8_sum + score_8_x608;
      res_9_sum <= res_9_sum + score_9_x608;
   end
   else if(res_done_x609) begin
      res_0_sum <= res_0_sum + score_0_x609;
      res_1_sum <= res_1_sum + score_1_x609;
      res_2_sum <= res_2_sum + score_2_x609;
      res_3_sum <= res_3_sum + score_3_x609;
      res_4_sum <= res_4_sum + score_4_x609;
      res_5_sum <= res_5_sum + score_5_x609;
      res_6_sum <= res_6_sum + score_6_x609;
      res_7_sum <= res_7_sum + score_7_x609;
      res_8_sum <= res_8_sum + score_8_x609;
      res_9_sum <= res_9_sum + score_9_x609;
   end
   else if(res_done_x610) begin
      res_0_sum <= res_0_sum + score_0_x610;
      res_1_sum <= res_1_sum + score_1_x610;
      res_2_sum <= res_2_sum + score_2_x610;
      res_3_sum <= res_3_sum + score_3_x610;
      res_4_sum <= res_4_sum + score_4_x610;
      res_5_sum <= res_5_sum + score_5_x610;
      res_6_sum <= res_6_sum + score_6_x610;
      res_7_sum <= res_7_sum + score_7_x610;
      res_8_sum <= res_8_sum + score_8_x610;
      res_9_sum <= res_9_sum + score_9_x610;
   end
   else if(res_done_x611) begin
      res_0_sum <= res_0_sum + score_0_x611;
      res_1_sum <= res_1_sum + score_1_x611;
      res_2_sum <= res_2_sum + score_2_x611;
      res_3_sum <= res_3_sum + score_3_x611;
      res_4_sum <= res_4_sum + score_4_x611;
      res_5_sum <= res_5_sum + score_5_x611;
      res_6_sum <= res_6_sum + score_6_x611;
      res_7_sum <= res_7_sum + score_7_x611;
      res_8_sum <= res_8_sum + score_8_x611;
      res_9_sum <= res_9_sum + score_9_x611;
   end
   else if(res_done_x612) begin
      res_0_sum <= res_0_sum + score_0_x612;
      res_1_sum <= res_1_sum + score_1_x612;
      res_2_sum <= res_2_sum + score_2_x612;
      res_3_sum <= res_3_sum + score_3_x612;
      res_4_sum <= res_4_sum + score_4_x612;
      res_5_sum <= res_5_sum + score_5_x612;
      res_6_sum <= res_6_sum + score_6_x612;
      res_7_sum <= res_7_sum + score_7_x612;
      res_8_sum <= res_8_sum + score_8_x612;
      res_9_sum <= res_9_sum + score_9_x612;
   end
   else if(res_done_x613) begin
      res_0_sum <= res_0_sum + score_0_x613;
      res_1_sum <= res_1_sum + score_1_x613;
      res_2_sum <= res_2_sum + score_2_x613;
      res_3_sum <= res_3_sum + score_3_x613;
      res_4_sum <= res_4_sum + score_4_x613;
      res_5_sum <= res_5_sum + score_5_x613;
      res_6_sum <= res_6_sum + score_6_x613;
      res_7_sum <= res_7_sum + score_7_x613;
      res_8_sum <= res_8_sum + score_8_x613;
      res_9_sum <= res_9_sum + score_9_x613;
   end
   else if(res_done_x614) begin
      res_0_sum <= res_0_sum + score_0_x614;
      res_1_sum <= res_1_sum + score_1_x614;
      res_2_sum <= res_2_sum + score_2_x614;
      res_3_sum <= res_3_sum + score_3_x614;
      res_4_sum <= res_4_sum + score_4_x614;
      res_5_sum <= res_5_sum + score_5_x614;
      res_6_sum <= res_6_sum + score_6_x614;
      res_7_sum <= res_7_sum + score_7_x614;
      res_8_sum <= res_8_sum + score_8_x614;
      res_9_sum <= res_9_sum + score_9_x614;
   end
   else if(res_done_x615) begin
      res_0_sum <= res_0_sum + score_0_x615;
      res_1_sum <= res_1_sum + score_1_x615;
      res_2_sum <= res_2_sum + score_2_x615;
      res_3_sum <= res_3_sum + score_3_x615;
      res_4_sum <= res_4_sum + score_4_x615;
      res_5_sum <= res_5_sum + score_5_x615;
      res_6_sum <= res_6_sum + score_6_x615;
      res_7_sum <= res_7_sum + score_7_x615;
      res_8_sum <= res_8_sum + score_8_x615;
      res_9_sum <= res_9_sum + score_9_x615;
   end
   else if(res_done_x616) begin
      res_0_sum <= res_0_sum + score_0_x616;
      res_1_sum <= res_1_sum + score_1_x616;
      res_2_sum <= res_2_sum + score_2_x616;
      res_3_sum <= res_3_sum + score_3_x616;
      res_4_sum <= res_4_sum + score_4_x616;
      res_5_sum <= res_5_sum + score_5_x616;
      res_6_sum <= res_6_sum + score_6_x616;
      res_7_sum <= res_7_sum + score_7_x616;
      res_8_sum <= res_8_sum + score_8_x616;
      res_9_sum <= res_9_sum + score_9_x616;
   end
   else if(res_done_x617) begin
      res_0_sum <= res_0_sum + score_0_x617;
      res_1_sum <= res_1_sum + score_1_x617;
      res_2_sum <= res_2_sum + score_2_x617;
      res_3_sum <= res_3_sum + score_3_x617;
      res_4_sum <= res_4_sum + score_4_x617;
      res_5_sum <= res_5_sum + score_5_x617;
      res_6_sum <= res_6_sum + score_6_x617;
      res_7_sum <= res_7_sum + score_7_x617;
      res_8_sum <= res_8_sum + score_8_x617;
      res_9_sum <= res_9_sum + score_9_x617;
   end
   else if(res_done_x618) begin
      res_0_sum <= res_0_sum + score_0_x618;
      res_1_sum <= res_1_sum + score_1_x618;
      res_2_sum <= res_2_sum + score_2_x618;
      res_3_sum <= res_3_sum + score_3_x618;
      res_4_sum <= res_4_sum + score_4_x618;
      res_5_sum <= res_5_sum + score_5_x618;
      res_6_sum <= res_6_sum + score_6_x618;
      res_7_sum <= res_7_sum + score_7_x618;
      res_8_sum <= res_8_sum + score_8_x618;
      res_9_sum <= res_9_sum + score_9_x618;
   end
   else if(res_done_x619) begin
      res_0_sum <= res_0_sum + score_0_x619;
      res_1_sum <= res_1_sum + score_1_x619;
      res_2_sum <= res_2_sum + score_2_x619;
      res_3_sum <= res_3_sum + score_3_x619;
      res_4_sum <= res_4_sum + score_4_x619;
      res_5_sum <= res_5_sum + score_5_x619;
      res_6_sum <= res_6_sum + score_6_x619;
      res_7_sum <= res_7_sum + score_7_x619;
      res_8_sum <= res_8_sum + score_8_x619;
      res_9_sum <= res_9_sum + score_9_x619;
   end
   else if(res_done_x620) begin
      res_0_sum <= res_0_sum + score_0_x620;
      res_1_sum <= res_1_sum + score_1_x620;
      res_2_sum <= res_2_sum + score_2_x620;
      res_3_sum <= res_3_sum + score_3_x620;
      res_4_sum <= res_4_sum + score_4_x620;
      res_5_sum <= res_5_sum + score_5_x620;
      res_6_sum <= res_6_sum + score_6_x620;
      res_7_sum <= res_7_sum + score_7_x620;
      res_8_sum <= res_8_sum + score_8_x620;
      res_9_sum <= res_9_sum + score_9_x620;
   end
   else if(res_done_x621) begin
      res_0_sum <= res_0_sum + score_0_x621;
      res_1_sum <= res_1_sum + score_1_x621;
      res_2_sum <= res_2_sum + score_2_x621;
      res_3_sum <= res_3_sum + score_3_x621;
      res_4_sum <= res_4_sum + score_4_x621;
      res_5_sum <= res_5_sum + score_5_x621;
      res_6_sum <= res_6_sum + score_6_x621;
      res_7_sum <= res_7_sum + score_7_x621;
      res_8_sum <= res_8_sum + score_8_x621;
      res_9_sum <= res_9_sum + score_9_x621;
   end
   else if(res_done_x622) begin
      res_0_sum <= res_0_sum + score_0_x622;
      res_1_sum <= res_1_sum + score_1_x622;
      res_2_sum <= res_2_sum + score_2_x622;
      res_3_sum <= res_3_sum + score_3_x622;
      res_4_sum <= res_4_sum + score_4_x622;
      res_5_sum <= res_5_sum + score_5_x622;
      res_6_sum <= res_6_sum + score_6_x622;
      res_7_sum <= res_7_sum + score_7_x622;
      res_8_sum <= res_8_sum + score_8_x622;
      res_9_sum <= res_9_sum + score_9_x622;
   end
   else if(res_done_x623) begin
      res_0_sum <= res_0_sum + score_0_x623;
      res_1_sum <= res_1_sum + score_1_x623;
      res_2_sum <= res_2_sum + score_2_x623;
      res_3_sum <= res_3_sum + score_3_x623;
      res_4_sum <= res_4_sum + score_4_x623;
      res_5_sum <= res_5_sum + score_5_x623;
      res_6_sum <= res_6_sum + score_6_x623;
      res_7_sum <= res_7_sum + score_7_x623;
      res_8_sum <= res_8_sum + score_8_x623;
      res_9_sum <= res_9_sum + score_9_x623;
   end
   else if(res_done_x624) begin
      res_0_sum <= res_0_sum + score_0_x624;
      res_1_sum <= res_1_sum + score_1_x624;
      res_2_sum <= res_2_sum + score_2_x624;
      res_3_sum <= res_3_sum + score_3_x624;
      res_4_sum <= res_4_sum + score_4_x624;
      res_5_sum <= res_5_sum + score_5_x624;
      res_6_sum <= res_6_sum + score_6_x624;
      res_7_sum <= res_7_sum + score_7_x624;
      res_8_sum <= res_8_sum + score_8_x624;
      res_9_sum <= res_9_sum + score_9_x624;
   end
   else if(res_done_x625) begin
      res_0_sum <= res_0_sum + score_0_x625;
      res_1_sum <= res_1_sum + score_1_x625;
      res_2_sum <= res_2_sum + score_2_x625;
      res_3_sum <= res_3_sum + score_3_x625;
      res_4_sum <= res_4_sum + score_4_x625;
      res_5_sum <= res_5_sum + score_5_x625;
      res_6_sum <= res_6_sum + score_6_x625;
      res_7_sum <= res_7_sum + score_7_x625;
      res_8_sum <= res_8_sum + score_8_x625;
      res_9_sum <= res_9_sum + score_9_x625;
   end
   else if(res_done_x626) begin
      res_0_sum <= res_0_sum + score_0_x626;
      res_1_sum <= res_1_sum + score_1_x626;
      res_2_sum <= res_2_sum + score_2_x626;
      res_3_sum <= res_3_sum + score_3_x626;
      res_4_sum <= res_4_sum + score_4_x626;
      res_5_sum <= res_5_sum + score_5_x626;
      res_6_sum <= res_6_sum + score_6_x626;
      res_7_sum <= res_7_sum + score_7_x626;
      res_8_sum <= res_8_sum + score_8_x626;
      res_9_sum <= res_9_sum + score_9_x626;
   end
   else if(res_done_x627) begin
      res_0_sum <= res_0_sum + score_0_x627;
      res_1_sum <= res_1_sum + score_1_x627;
      res_2_sum <= res_2_sum + score_2_x627;
      res_3_sum <= res_3_sum + score_3_x627;
      res_4_sum <= res_4_sum + score_4_x627;
      res_5_sum <= res_5_sum + score_5_x627;
      res_6_sum <= res_6_sum + score_6_x627;
      res_7_sum <= res_7_sum + score_7_x627;
      res_8_sum <= res_8_sum + score_8_x627;
      res_9_sum <= res_9_sum + score_9_x627;
   end
   else if(res_done_x628) begin
      res_0_sum <= res_0_sum + score_0_x628;
      res_1_sum <= res_1_sum + score_1_x628;
      res_2_sum <= res_2_sum + score_2_x628;
      res_3_sum <= res_3_sum + score_3_x628;
      res_4_sum <= res_4_sum + score_4_x628;
      res_5_sum <= res_5_sum + score_5_x628;
      res_6_sum <= res_6_sum + score_6_x628;
      res_7_sum <= res_7_sum + score_7_x628;
      res_8_sum <= res_8_sum + score_8_x628;
      res_9_sum <= res_9_sum + score_9_x628;
   end
   else if(res_done_x629) begin
      res_0_sum <= res_0_sum + score_0_x629;
      res_1_sum <= res_1_sum + score_1_x629;
      res_2_sum <= res_2_sum + score_2_x629;
      res_3_sum <= res_3_sum + score_3_x629;
      res_4_sum <= res_4_sum + score_4_x629;
      res_5_sum <= res_5_sum + score_5_x629;
      res_6_sum <= res_6_sum + score_6_x629;
      res_7_sum <= res_7_sum + score_7_x629;
      res_8_sum <= res_8_sum + score_8_x629;
      res_9_sum <= res_9_sum + score_9_x629;
   end
   else if(res_done_x630) begin
      res_0_sum <= res_0_sum + score_0_x630;
      res_1_sum <= res_1_sum + score_1_x630;
      res_2_sum <= res_2_sum + score_2_x630;
      res_3_sum <= res_3_sum + score_3_x630;
      res_4_sum <= res_4_sum + score_4_x630;
      res_5_sum <= res_5_sum + score_5_x630;
      res_6_sum <= res_6_sum + score_6_x630;
      res_7_sum <= res_7_sum + score_7_x630;
      res_8_sum <= res_8_sum + score_8_x630;
      res_9_sum <= res_9_sum + score_9_x630;
   end
   else if(res_done_x631) begin
      res_0_sum <= res_0_sum + score_0_x631;
      res_1_sum <= res_1_sum + score_1_x631;
      res_2_sum <= res_2_sum + score_2_x631;
      res_3_sum <= res_3_sum + score_3_x631;
      res_4_sum <= res_4_sum + score_4_x631;
      res_5_sum <= res_5_sum + score_5_x631;
      res_6_sum <= res_6_sum + score_6_x631;
      res_7_sum <= res_7_sum + score_7_x631;
      res_8_sum <= res_8_sum + score_8_x631;
      res_9_sum <= res_9_sum + score_9_x631;
   end
   else if(res_done_x632) begin
      res_0_sum <= res_0_sum + score_0_x632;
      res_1_sum <= res_1_sum + score_1_x632;
      res_2_sum <= res_2_sum + score_2_x632;
      res_3_sum <= res_3_sum + score_3_x632;
      res_4_sum <= res_4_sum + score_4_x632;
      res_5_sum <= res_5_sum + score_5_x632;
      res_6_sum <= res_6_sum + score_6_x632;
      res_7_sum <= res_7_sum + score_7_x632;
      res_8_sum <= res_8_sum + score_8_x632;
      res_9_sum <= res_9_sum + score_9_x632;
   end
   else if(res_done_x633) begin
      res_0_sum <= res_0_sum + score_0_x633;
      res_1_sum <= res_1_sum + score_1_x633;
      res_2_sum <= res_2_sum + score_2_x633;
      res_3_sum <= res_3_sum + score_3_x633;
      res_4_sum <= res_4_sum + score_4_x633;
      res_5_sum <= res_5_sum + score_5_x633;
      res_6_sum <= res_6_sum + score_6_x633;
      res_7_sum <= res_7_sum + score_7_x633;
      res_8_sum <= res_8_sum + score_8_x633;
      res_9_sum <= res_9_sum + score_9_x633;
   end
   else if(res_done_x634) begin
      res_0_sum <= res_0_sum + score_0_x634;
      res_1_sum <= res_1_sum + score_1_x634;
      res_2_sum <= res_2_sum + score_2_x634;
      res_3_sum <= res_3_sum + score_3_x634;
      res_4_sum <= res_4_sum + score_4_x634;
      res_5_sum <= res_5_sum + score_5_x634;
      res_6_sum <= res_6_sum + score_6_x634;
      res_7_sum <= res_7_sum + score_7_x634;
      res_8_sum <= res_8_sum + score_8_x634;
      res_9_sum <= res_9_sum + score_9_x634;
   end
   else if(res_done_x635) begin
      res_0_sum <= res_0_sum + score_0_x635;
      res_1_sum <= res_1_sum + score_1_x635;
      res_2_sum <= res_2_sum + score_2_x635;
      res_3_sum <= res_3_sum + score_3_x635;
      res_4_sum <= res_4_sum + score_4_x635;
      res_5_sum <= res_5_sum + score_5_x635;
      res_6_sum <= res_6_sum + score_6_x635;
      res_7_sum <= res_7_sum + score_7_x635;
      res_8_sum <= res_8_sum + score_8_x635;
      res_9_sum <= res_9_sum + score_9_x635;
   end
   else if(res_done_x636) begin
      res_0_sum <= res_0_sum + score_0_x636;
      res_1_sum <= res_1_sum + score_1_x636;
      res_2_sum <= res_2_sum + score_2_x636;
      res_3_sum <= res_3_sum + score_3_x636;
      res_4_sum <= res_4_sum + score_4_x636;
      res_5_sum <= res_5_sum + score_5_x636;
      res_6_sum <= res_6_sum + score_6_x636;
      res_7_sum <= res_7_sum + score_7_x636;
      res_8_sum <= res_8_sum + score_8_x636;
      res_9_sum <= res_9_sum + score_9_x636;
   end
   else if(res_done_x637) begin
      res_0_sum <= res_0_sum + score_0_x637;
      res_1_sum <= res_1_sum + score_1_x637;
      res_2_sum <= res_2_sum + score_2_x637;
      res_3_sum <= res_3_sum + score_3_x637;
      res_4_sum <= res_4_sum + score_4_x637;
      res_5_sum <= res_5_sum + score_5_x637;
      res_6_sum <= res_6_sum + score_6_x637;
      res_7_sum <= res_7_sum + score_7_x637;
      res_8_sum <= res_8_sum + score_8_x637;
      res_9_sum <= res_9_sum + score_9_x637;
   end
   else if(res_done_x638) begin
      res_0_sum <= res_0_sum + score_0_x638;
      res_1_sum <= res_1_sum + score_1_x638;
      res_2_sum <= res_2_sum + score_2_x638;
      res_3_sum <= res_3_sum + score_3_x638;
      res_4_sum <= res_4_sum + score_4_x638;
      res_5_sum <= res_5_sum + score_5_x638;
      res_6_sum <= res_6_sum + score_6_x638;
      res_7_sum <= res_7_sum + score_7_x638;
      res_8_sum <= res_8_sum + score_8_x638;
      res_9_sum <= res_9_sum + score_9_x638;
   end
   else if(res_done_x639) begin
      res_0_sum <= res_0_sum + score_0_x639;
      res_1_sum <= res_1_sum + score_1_x639;
      res_2_sum <= res_2_sum + score_2_x639;
      res_3_sum <= res_3_sum + score_3_x639;
      res_4_sum <= res_4_sum + score_4_x639;
      res_5_sum <= res_5_sum + score_5_x639;
      res_6_sum <= res_6_sum + score_6_x639;
      res_7_sum <= res_7_sum + score_7_x639;
      res_8_sum <= res_8_sum + score_8_x639;
      res_9_sum <= res_9_sum + score_9_x639;
   end
   else if(res_done_x640) begin
      res_0_sum <= res_0_sum + score_0_x640;
      res_1_sum <= res_1_sum + score_1_x640;
      res_2_sum <= res_2_sum + score_2_x640;
      res_3_sum <= res_3_sum + score_3_x640;
      res_4_sum <= res_4_sum + score_4_x640;
      res_5_sum <= res_5_sum + score_5_x640;
      res_6_sum <= res_6_sum + score_6_x640;
      res_7_sum <= res_7_sum + score_7_x640;
      res_8_sum <= res_8_sum + score_8_x640;
      res_9_sum <= res_9_sum + score_9_x640;
   end
   else if(res_done_x641) begin
      res_0_sum <= res_0_sum + score_0_x641;
      res_1_sum <= res_1_sum + score_1_x641;
      res_2_sum <= res_2_sum + score_2_x641;
      res_3_sum <= res_3_sum + score_3_x641;
      res_4_sum <= res_4_sum + score_4_x641;
      res_5_sum <= res_5_sum + score_5_x641;
      res_6_sum <= res_6_sum + score_6_x641;
      res_7_sum <= res_7_sum + score_7_x641;
      res_8_sum <= res_8_sum + score_8_x641;
      res_9_sum <= res_9_sum + score_9_x641;
   end
   else if(res_done_x642) begin
      res_0_sum <= res_0_sum + score_0_x642;
      res_1_sum <= res_1_sum + score_1_x642;
      res_2_sum <= res_2_sum + score_2_x642;
      res_3_sum <= res_3_sum + score_3_x642;
      res_4_sum <= res_4_sum + score_4_x642;
      res_5_sum <= res_5_sum + score_5_x642;
      res_6_sum <= res_6_sum + score_6_x642;
      res_7_sum <= res_7_sum + score_7_x642;
      res_8_sum <= res_8_sum + score_8_x642;
      res_9_sum <= res_9_sum + score_9_x642;
   end
   else if(res_done_x643) begin
      res_0_sum <= res_0_sum + score_0_x643;
      res_1_sum <= res_1_sum + score_1_x643;
      res_2_sum <= res_2_sum + score_2_x643;
      res_3_sum <= res_3_sum + score_3_x643;
      res_4_sum <= res_4_sum + score_4_x643;
      res_5_sum <= res_5_sum + score_5_x643;
      res_6_sum <= res_6_sum + score_6_x643;
      res_7_sum <= res_7_sum + score_7_x643;
      res_8_sum <= res_8_sum + score_8_x643;
      res_9_sum <= res_9_sum + score_9_x643;
   end
   else if(res_done_x644) begin
      res_0_sum <= res_0_sum + score_0_x644;
      res_1_sum <= res_1_sum + score_1_x644;
      res_2_sum <= res_2_sum + score_2_x644;
      res_3_sum <= res_3_sum + score_3_x644;
      res_4_sum <= res_4_sum + score_4_x644;
      res_5_sum <= res_5_sum + score_5_x644;
      res_6_sum <= res_6_sum + score_6_x644;
      res_7_sum <= res_7_sum + score_7_x644;
      res_8_sum <= res_8_sum + score_8_x644;
      res_9_sum <= res_9_sum + score_9_x644;
   end
   else if(res_done_x645) begin
      res_0_sum <= res_0_sum + score_0_x645;
      res_1_sum <= res_1_sum + score_1_x645;
      res_2_sum <= res_2_sum + score_2_x645;
      res_3_sum <= res_3_sum + score_3_x645;
      res_4_sum <= res_4_sum + score_4_x645;
      res_5_sum <= res_5_sum + score_5_x645;
      res_6_sum <= res_6_sum + score_6_x645;
      res_7_sum <= res_7_sum + score_7_x645;
      res_8_sum <= res_8_sum + score_8_x645;
      res_9_sum <= res_9_sum + score_9_x645;
   end
   else if(res_done_x646) begin
      res_0_sum <= res_0_sum + score_0_x646;
      res_1_sum <= res_1_sum + score_1_x646;
      res_2_sum <= res_2_sum + score_2_x646;
      res_3_sum <= res_3_sum + score_3_x646;
      res_4_sum <= res_4_sum + score_4_x646;
      res_5_sum <= res_5_sum + score_5_x646;
      res_6_sum <= res_6_sum + score_6_x646;
      res_7_sum <= res_7_sum + score_7_x646;
      res_8_sum <= res_8_sum + score_8_x646;
      res_9_sum <= res_9_sum + score_9_x646;
   end
   else if(res_done_x647) begin
      res_0_sum <= res_0_sum + score_0_x647;
      res_1_sum <= res_1_sum + score_1_x647;
      res_2_sum <= res_2_sum + score_2_x647;
      res_3_sum <= res_3_sum + score_3_x647;
      res_4_sum <= res_4_sum + score_4_x647;
      res_5_sum <= res_5_sum + score_5_x647;
      res_6_sum <= res_6_sum + score_6_x647;
      res_7_sum <= res_7_sum + score_7_x647;
      res_8_sum <= res_8_sum + score_8_x647;
      res_9_sum <= res_9_sum + score_9_x647;
   end
   else if(res_done_x648) begin
      res_0_sum <= res_0_sum + score_0_x648;
      res_1_sum <= res_1_sum + score_1_x648;
      res_2_sum <= res_2_sum + score_2_x648;
      res_3_sum <= res_3_sum + score_3_x648;
      res_4_sum <= res_4_sum + score_4_x648;
      res_5_sum <= res_5_sum + score_5_x648;
      res_6_sum <= res_6_sum + score_6_x648;
      res_7_sum <= res_7_sum + score_7_x648;
      res_8_sum <= res_8_sum + score_8_x648;
      res_9_sum <= res_9_sum + score_9_x648;
   end
   else if(res_done_x649) begin
      res_0_sum <= res_0_sum + score_0_x649;
      res_1_sum <= res_1_sum + score_1_x649;
      res_2_sum <= res_2_sum + score_2_x649;
      res_3_sum <= res_3_sum + score_3_x649;
      res_4_sum <= res_4_sum + score_4_x649;
      res_5_sum <= res_5_sum + score_5_x649;
      res_6_sum <= res_6_sum + score_6_x649;
      res_7_sum <= res_7_sum + score_7_x649;
      res_8_sum <= res_8_sum + score_8_x649;
      res_9_sum <= res_9_sum + score_9_x649;
   end
   else if(res_done_x650) begin
      res_0_sum <= res_0_sum + score_0_x650;
      res_1_sum <= res_1_sum + score_1_x650;
      res_2_sum <= res_2_sum + score_2_x650;
      res_3_sum <= res_3_sum + score_3_x650;
      res_4_sum <= res_4_sum + score_4_x650;
      res_5_sum <= res_5_sum + score_5_x650;
      res_6_sum <= res_6_sum + score_6_x650;
      res_7_sum <= res_7_sum + score_7_x650;
      res_8_sum <= res_8_sum + score_8_x650;
      res_9_sum <= res_9_sum + score_9_x650;
   end
   else if(res_done_x651) begin
      res_0_sum <= res_0_sum + score_0_x651;
      res_1_sum <= res_1_sum + score_1_x651;
      res_2_sum <= res_2_sum + score_2_x651;
      res_3_sum <= res_3_sum + score_3_x651;
      res_4_sum <= res_4_sum + score_4_x651;
      res_5_sum <= res_5_sum + score_5_x651;
      res_6_sum <= res_6_sum + score_6_x651;
      res_7_sum <= res_7_sum + score_7_x651;
      res_8_sum <= res_8_sum + score_8_x651;
      res_9_sum <= res_9_sum + score_9_x651;
   end
   else if(res_done_x652) begin
      res_0_sum <= res_0_sum + score_0_x652;
      res_1_sum <= res_1_sum + score_1_x652;
      res_2_sum <= res_2_sum + score_2_x652;
      res_3_sum <= res_3_sum + score_3_x652;
      res_4_sum <= res_4_sum + score_4_x652;
      res_5_sum <= res_5_sum + score_5_x652;
      res_6_sum <= res_6_sum + score_6_x652;
      res_7_sum <= res_7_sum + score_7_x652;
      res_8_sum <= res_8_sum + score_8_x652;
      res_9_sum <= res_9_sum + score_9_x652;
   end
   else if(res_done_x653) begin
      res_0_sum <= res_0_sum + score_0_x653;
      res_1_sum <= res_1_sum + score_1_x653;
      res_2_sum <= res_2_sum + score_2_x653;
      res_3_sum <= res_3_sum + score_3_x653;
      res_4_sum <= res_4_sum + score_4_x653;
      res_5_sum <= res_5_sum + score_5_x653;
      res_6_sum <= res_6_sum + score_6_x653;
      res_7_sum <= res_7_sum + score_7_x653;
      res_8_sum <= res_8_sum + score_8_x653;
      res_9_sum <= res_9_sum + score_9_x653;
   end
   else if(res_done_x654) begin
      res_0_sum <= res_0_sum + score_0_x654;
      res_1_sum <= res_1_sum + score_1_x654;
      res_2_sum <= res_2_sum + score_2_x654;
      res_3_sum <= res_3_sum + score_3_x654;
      res_4_sum <= res_4_sum + score_4_x654;
      res_5_sum <= res_5_sum + score_5_x654;
      res_6_sum <= res_6_sum + score_6_x654;
      res_7_sum <= res_7_sum + score_7_x654;
      res_8_sum <= res_8_sum + score_8_x654;
      res_9_sum <= res_9_sum + score_9_x654;
   end
   else if(res_done_x655) begin
      res_0_sum <= res_0_sum + score_0_x655;
      res_1_sum <= res_1_sum + score_1_x655;
      res_2_sum <= res_2_sum + score_2_x655;
      res_3_sum <= res_3_sum + score_3_x655;
      res_4_sum <= res_4_sum + score_4_x655;
      res_5_sum <= res_5_sum + score_5_x655;
      res_6_sum <= res_6_sum + score_6_x655;
      res_7_sum <= res_7_sum + score_7_x655;
      res_8_sum <= res_8_sum + score_8_x655;
      res_9_sum <= res_9_sum + score_9_x655;
   end
   else if(res_done_x656) begin
      res_0_sum <= res_0_sum + score_0_x656;
      res_1_sum <= res_1_sum + score_1_x656;
      res_2_sum <= res_2_sum + score_2_x656;
      res_3_sum <= res_3_sum + score_3_x656;
      res_4_sum <= res_4_sum + score_4_x656;
      res_5_sum <= res_5_sum + score_5_x656;
      res_6_sum <= res_6_sum + score_6_x656;
      res_7_sum <= res_7_sum + score_7_x656;
      res_8_sum <= res_8_sum + score_8_x656;
      res_9_sum <= res_9_sum + score_9_x656;
   end
   else if(res_done_x657) begin
      res_0_sum <= res_0_sum + score_0_x657;
      res_1_sum <= res_1_sum + score_1_x657;
      res_2_sum <= res_2_sum + score_2_x657;
      res_3_sum <= res_3_sum + score_3_x657;
      res_4_sum <= res_4_sum + score_4_x657;
      res_5_sum <= res_5_sum + score_5_x657;
      res_6_sum <= res_6_sum + score_6_x657;
      res_7_sum <= res_7_sum + score_7_x657;
      res_8_sum <= res_8_sum + score_8_x657;
      res_9_sum <= res_9_sum + score_9_x657;
   end
   else if(res_done_x658) begin
      res_0_sum <= res_0_sum + score_0_x658;
      res_1_sum <= res_1_sum + score_1_x658;
      res_2_sum <= res_2_sum + score_2_x658;
      res_3_sum <= res_3_sum + score_3_x658;
      res_4_sum <= res_4_sum + score_4_x658;
      res_5_sum <= res_5_sum + score_5_x658;
      res_6_sum <= res_6_sum + score_6_x658;
      res_7_sum <= res_7_sum + score_7_x658;
      res_8_sum <= res_8_sum + score_8_x658;
      res_9_sum <= res_9_sum + score_9_x658;
   end
   else if(res_done_x659) begin
      res_0_sum <= res_0_sum + score_0_x659;
      res_1_sum <= res_1_sum + score_1_x659;
      res_2_sum <= res_2_sum + score_2_x659;
      res_3_sum <= res_3_sum + score_3_x659;
      res_4_sum <= res_4_sum + score_4_x659;
      res_5_sum <= res_5_sum + score_5_x659;
      res_6_sum <= res_6_sum + score_6_x659;
      res_7_sum <= res_7_sum + score_7_x659;
      res_8_sum <= res_8_sum + score_8_x659;
      res_9_sum <= res_9_sum + score_9_x659;
   end
   else if(res_done_x660) begin
      res_0_sum <= res_0_sum + score_0_x660;
      res_1_sum <= res_1_sum + score_1_x660;
      res_2_sum <= res_2_sum + score_2_x660;
      res_3_sum <= res_3_sum + score_3_x660;
      res_4_sum <= res_4_sum + score_4_x660;
      res_5_sum <= res_5_sum + score_5_x660;
      res_6_sum <= res_6_sum + score_6_x660;
      res_7_sum <= res_7_sum + score_7_x660;
      res_8_sum <= res_8_sum + score_8_x660;
      res_9_sum <= res_9_sum + score_9_x660;
   end
   else if(res_done_x661) begin
      res_0_sum <= res_0_sum + score_0_x661;
      res_1_sum <= res_1_sum + score_1_x661;
      res_2_sum <= res_2_sum + score_2_x661;
      res_3_sum <= res_3_sum + score_3_x661;
      res_4_sum <= res_4_sum + score_4_x661;
      res_5_sum <= res_5_sum + score_5_x661;
      res_6_sum <= res_6_sum + score_6_x661;
      res_7_sum <= res_7_sum + score_7_x661;
      res_8_sum <= res_8_sum + score_8_x661;
      res_9_sum <= res_9_sum + score_9_x661;
   end
   else if(res_done_x662) begin
      res_0_sum <= res_0_sum + score_0_x662;
      res_1_sum <= res_1_sum + score_1_x662;
      res_2_sum <= res_2_sum + score_2_x662;
      res_3_sum <= res_3_sum + score_3_x662;
      res_4_sum <= res_4_sum + score_4_x662;
      res_5_sum <= res_5_sum + score_5_x662;
      res_6_sum <= res_6_sum + score_6_x662;
      res_7_sum <= res_7_sum + score_7_x662;
      res_8_sum <= res_8_sum + score_8_x662;
      res_9_sum <= res_9_sum + score_9_x662;
   end
   else if(res_done_x663) begin
      res_0_sum <= res_0_sum + score_0_x663;
      res_1_sum <= res_1_sum + score_1_x663;
      res_2_sum <= res_2_sum + score_2_x663;
      res_3_sum <= res_3_sum + score_3_x663;
      res_4_sum <= res_4_sum + score_4_x663;
      res_5_sum <= res_5_sum + score_5_x663;
      res_6_sum <= res_6_sum + score_6_x663;
      res_7_sum <= res_7_sum + score_7_x663;
      res_8_sum <= res_8_sum + score_8_x663;
      res_9_sum <= res_9_sum + score_9_x663;
   end
   else if(res_done_x664) begin
      res_0_sum <= res_0_sum + score_0_x664;
      res_1_sum <= res_1_sum + score_1_x664;
      res_2_sum <= res_2_sum + score_2_x664;
      res_3_sum <= res_3_sum + score_3_x664;
      res_4_sum <= res_4_sum + score_4_x664;
      res_5_sum <= res_5_sum + score_5_x664;
      res_6_sum <= res_6_sum + score_6_x664;
      res_7_sum <= res_7_sum + score_7_x664;
      res_8_sum <= res_8_sum + score_8_x664;
      res_9_sum <= res_9_sum + score_9_x664;
   end
   else if(res_done_x665) begin
      res_0_sum <= res_0_sum + score_0_x665;
      res_1_sum <= res_1_sum + score_1_x665;
      res_2_sum <= res_2_sum + score_2_x665;
      res_3_sum <= res_3_sum + score_3_x665;
      res_4_sum <= res_4_sum + score_4_x665;
      res_5_sum <= res_5_sum + score_5_x665;
      res_6_sum <= res_6_sum + score_6_x665;
      res_7_sum <= res_7_sum + score_7_x665;
      res_8_sum <= res_8_sum + score_8_x665;
      res_9_sum <= res_9_sum + score_9_x665;
   end
   else if(res_done_x666) begin
      res_0_sum <= res_0_sum + score_0_x666;
      res_1_sum <= res_1_sum + score_1_x666;
      res_2_sum <= res_2_sum + score_2_x666;
      res_3_sum <= res_3_sum + score_3_x666;
      res_4_sum <= res_4_sum + score_4_x666;
      res_5_sum <= res_5_sum + score_5_x666;
      res_6_sum <= res_6_sum + score_6_x666;
      res_7_sum <= res_7_sum + score_7_x666;
      res_8_sum <= res_8_sum + score_8_x666;
      res_9_sum <= res_9_sum + score_9_x666;
   end
   else if(res_done_x667) begin
      res_0_sum <= res_0_sum + score_0_x667;
      res_1_sum <= res_1_sum + score_1_x667;
      res_2_sum <= res_2_sum + score_2_x667;
      res_3_sum <= res_3_sum + score_3_x667;
      res_4_sum <= res_4_sum + score_4_x667;
      res_5_sum <= res_5_sum + score_5_x667;
      res_6_sum <= res_6_sum + score_6_x667;
      res_7_sum <= res_7_sum + score_7_x667;
      res_8_sum <= res_8_sum + score_8_x667;
      res_9_sum <= res_9_sum + score_9_x667;
   end
   else if(res_done_x668) begin
      res_0_sum <= res_0_sum + score_0_x668;
      res_1_sum <= res_1_sum + score_1_x668;
      res_2_sum <= res_2_sum + score_2_x668;
      res_3_sum <= res_3_sum + score_3_x668;
      res_4_sum <= res_4_sum + score_4_x668;
      res_5_sum <= res_5_sum + score_5_x668;
      res_6_sum <= res_6_sum + score_6_x668;
      res_7_sum <= res_7_sum + score_7_x668;
      res_8_sum <= res_8_sum + score_8_x668;
      res_9_sum <= res_9_sum + score_9_x668;
   end
   else if(res_done_x669) begin
      res_0_sum <= res_0_sum + score_0_x669;
      res_1_sum <= res_1_sum + score_1_x669;
      res_2_sum <= res_2_sum + score_2_x669;
      res_3_sum <= res_3_sum + score_3_x669;
      res_4_sum <= res_4_sum + score_4_x669;
      res_5_sum <= res_5_sum + score_5_x669;
      res_6_sum <= res_6_sum + score_6_x669;
      res_7_sum <= res_7_sum + score_7_x669;
      res_8_sum <= res_8_sum + score_8_x669;
      res_9_sum <= res_9_sum + score_9_x669;
   end
   else if(res_done_x670) begin
      res_0_sum <= res_0_sum + score_0_x670;
      res_1_sum <= res_1_sum + score_1_x670;
      res_2_sum <= res_2_sum + score_2_x670;
      res_3_sum <= res_3_sum + score_3_x670;
      res_4_sum <= res_4_sum + score_4_x670;
      res_5_sum <= res_5_sum + score_5_x670;
      res_6_sum <= res_6_sum + score_6_x670;
      res_7_sum <= res_7_sum + score_7_x670;
      res_8_sum <= res_8_sum + score_8_x670;
      res_9_sum <= res_9_sum + score_9_x670;
   end
   else if(res_done_x671) begin
      res_0_sum <= res_0_sum + score_0_x671;
      res_1_sum <= res_1_sum + score_1_x671;
      res_2_sum <= res_2_sum + score_2_x671;
      res_3_sum <= res_3_sum + score_3_x671;
      res_4_sum <= res_4_sum + score_4_x671;
      res_5_sum <= res_5_sum + score_5_x671;
      res_6_sum <= res_6_sum + score_6_x671;
      res_7_sum <= res_7_sum + score_7_x671;
      res_8_sum <= res_8_sum + score_8_x671;
      res_9_sum <= res_9_sum + score_9_x671;
   end
   else if(res_done_x672) begin
      res_0_sum <= res_0_sum + score_0_x672;
      res_1_sum <= res_1_sum + score_1_x672;
      res_2_sum <= res_2_sum + score_2_x672;
      res_3_sum <= res_3_sum + score_3_x672;
      res_4_sum <= res_4_sum + score_4_x672;
      res_5_sum <= res_5_sum + score_5_x672;
      res_6_sum <= res_6_sum + score_6_x672;
      res_7_sum <= res_7_sum + score_7_x672;
      res_8_sum <= res_8_sum + score_8_x672;
      res_9_sum <= res_9_sum + score_9_x672;
   end
   else if(res_done_x673) begin
      res_0_sum <= res_0_sum + score_0_x673;
      res_1_sum <= res_1_sum + score_1_x673;
      res_2_sum <= res_2_sum + score_2_x673;
      res_3_sum <= res_3_sum + score_3_x673;
      res_4_sum <= res_4_sum + score_4_x673;
      res_5_sum <= res_5_sum + score_5_x673;
      res_6_sum <= res_6_sum + score_6_x673;
      res_7_sum <= res_7_sum + score_7_x673;
      res_8_sum <= res_8_sum + score_8_x673;
      res_9_sum <= res_9_sum + score_9_x673;
   end
   else if(res_done_x674) begin
      res_0_sum <= res_0_sum + score_0_x674;
      res_1_sum <= res_1_sum + score_1_x674;
      res_2_sum <= res_2_sum + score_2_x674;
      res_3_sum <= res_3_sum + score_3_x674;
      res_4_sum <= res_4_sum + score_4_x674;
      res_5_sum <= res_5_sum + score_5_x674;
      res_6_sum <= res_6_sum + score_6_x674;
      res_7_sum <= res_7_sum + score_7_x674;
      res_8_sum <= res_8_sum + score_8_x674;
      res_9_sum <= res_9_sum + score_9_x674;
   end
   else if(res_done_x675) begin
      res_0_sum <= res_0_sum + score_0_x675;
      res_1_sum <= res_1_sum + score_1_x675;
      res_2_sum <= res_2_sum + score_2_x675;
      res_3_sum <= res_3_sum + score_3_x675;
      res_4_sum <= res_4_sum + score_4_x675;
      res_5_sum <= res_5_sum + score_5_x675;
      res_6_sum <= res_6_sum + score_6_x675;
      res_7_sum <= res_7_sum + score_7_x675;
      res_8_sum <= res_8_sum + score_8_x675;
      res_9_sum <= res_9_sum + score_9_x675;
   end
   else if(res_done_x676) begin
      res_0_sum <= res_0_sum + score_0_x676;
      res_1_sum <= res_1_sum + score_1_x676;
      res_2_sum <= res_2_sum + score_2_x676;
      res_3_sum <= res_3_sum + score_3_x676;
      res_4_sum <= res_4_sum + score_4_x676;
      res_5_sum <= res_5_sum + score_5_x676;
      res_6_sum <= res_6_sum + score_6_x676;
      res_7_sum <= res_7_sum + score_7_x676;
      res_8_sum <= res_8_sum + score_8_x676;
      res_9_sum <= res_9_sum + score_9_x676;
   end
   else if(res_done_x677) begin
      res_0_sum <= res_0_sum + score_0_x677;
      res_1_sum <= res_1_sum + score_1_x677;
      res_2_sum <= res_2_sum + score_2_x677;
      res_3_sum <= res_3_sum + score_3_x677;
      res_4_sum <= res_4_sum + score_4_x677;
      res_5_sum <= res_5_sum + score_5_x677;
      res_6_sum <= res_6_sum + score_6_x677;
      res_7_sum <= res_7_sum + score_7_x677;
      res_8_sum <= res_8_sum + score_8_x677;
      res_9_sum <= res_9_sum + score_9_x677;
   end
   else if(res_done_x678) begin
      res_0_sum <= res_0_sum + score_0_x678;
      res_1_sum <= res_1_sum + score_1_x678;
      res_2_sum <= res_2_sum + score_2_x678;
      res_3_sum <= res_3_sum + score_3_x678;
      res_4_sum <= res_4_sum + score_4_x678;
      res_5_sum <= res_5_sum + score_5_x678;
      res_6_sum <= res_6_sum + score_6_x678;
      res_7_sum <= res_7_sum + score_7_x678;
      res_8_sum <= res_8_sum + score_8_x678;
      res_9_sum <= res_9_sum + score_9_x678;
   end
   else if(res_done_x679) begin
      res_0_sum <= res_0_sum + score_0_x679;
      res_1_sum <= res_1_sum + score_1_x679;
      res_2_sum <= res_2_sum + score_2_x679;
      res_3_sum <= res_3_sum + score_3_x679;
      res_4_sum <= res_4_sum + score_4_x679;
      res_5_sum <= res_5_sum + score_5_x679;
      res_6_sum <= res_6_sum + score_6_x679;
      res_7_sum <= res_7_sum + score_7_x679;
      res_8_sum <= res_8_sum + score_8_x679;
      res_9_sum <= res_9_sum + score_9_x679;
   end
   else if(res_done_x680) begin
      res_0_sum <= res_0_sum + score_0_x680;
      res_1_sum <= res_1_sum + score_1_x680;
      res_2_sum <= res_2_sum + score_2_x680;
      res_3_sum <= res_3_sum + score_3_x680;
      res_4_sum <= res_4_sum + score_4_x680;
      res_5_sum <= res_5_sum + score_5_x680;
      res_6_sum <= res_6_sum + score_6_x680;
      res_7_sum <= res_7_sum + score_7_x680;
      res_8_sum <= res_8_sum + score_8_x680;
      res_9_sum <= res_9_sum + score_9_x680;
   end
   else if(res_done_x681) begin
      res_0_sum <= res_0_sum + score_0_x681;
      res_1_sum <= res_1_sum + score_1_x681;
      res_2_sum <= res_2_sum + score_2_x681;
      res_3_sum <= res_3_sum + score_3_x681;
      res_4_sum <= res_4_sum + score_4_x681;
      res_5_sum <= res_5_sum + score_5_x681;
      res_6_sum <= res_6_sum + score_6_x681;
      res_7_sum <= res_7_sum + score_7_x681;
      res_8_sum <= res_8_sum + score_8_x681;
      res_9_sum <= res_9_sum + score_9_x681;
   end
   else if(res_done_x682) begin
      res_0_sum <= res_0_sum + score_0_x682;
      res_1_sum <= res_1_sum + score_1_x682;
      res_2_sum <= res_2_sum + score_2_x682;
      res_3_sum <= res_3_sum + score_3_x682;
      res_4_sum <= res_4_sum + score_4_x682;
      res_5_sum <= res_5_sum + score_5_x682;
      res_6_sum <= res_6_sum + score_6_x682;
      res_7_sum <= res_7_sum + score_7_x682;
      res_8_sum <= res_8_sum + score_8_x682;
      res_9_sum <= res_9_sum + score_9_x682;
   end
   else if(res_done_x683) begin
      res_0_sum <= res_0_sum + score_0_x683;
      res_1_sum <= res_1_sum + score_1_x683;
      res_2_sum <= res_2_sum + score_2_x683;
      res_3_sum <= res_3_sum + score_3_x683;
      res_4_sum <= res_4_sum + score_4_x683;
      res_5_sum <= res_5_sum + score_5_x683;
      res_6_sum <= res_6_sum + score_6_x683;
      res_7_sum <= res_7_sum + score_7_x683;
      res_8_sum <= res_8_sum + score_8_x683;
      res_9_sum <= res_9_sum + score_9_x683;
   end
   else if(res_done_x684) begin
      res_0_sum <= res_0_sum + score_0_x684;
      res_1_sum <= res_1_sum + score_1_x684;
      res_2_sum <= res_2_sum + score_2_x684;
      res_3_sum <= res_3_sum + score_3_x684;
      res_4_sum <= res_4_sum + score_4_x684;
      res_5_sum <= res_5_sum + score_5_x684;
      res_6_sum <= res_6_sum + score_6_x684;
      res_7_sum <= res_7_sum + score_7_x684;
      res_8_sum <= res_8_sum + score_8_x684;
      res_9_sum <= res_9_sum + score_9_x684;
   end
   else if(res_done_x685) begin
      res_0_sum <= res_0_sum + score_0_x685;
      res_1_sum <= res_1_sum + score_1_x685;
      res_2_sum <= res_2_sum + score_2_x685;
      res_3_sum <= res_3_sum + score_3_x685;
      res_4_sum <= res_4_sum + score_4_x685;
      res_5_sum <= res_5_sum + score_5_x685;
      res_6_sum <= res_6_sum + score_6_x685;
      res_7_sum <= res_7_sum + score_7_x685;
      res_8_sum <= res_8_sum + score_8_x685;
      res_9_sum <= res_9_sum + score_9_x685;
   end
   else if(res_done_x686) begin
      res_0_sum <= res_0_sum + score_0_x686;
      res_1_sum <= res_1_sum + score_1_x686;
      res_2_sum <= res_2_sum + score_2_x686;
      res_3_sum <= res_3_sum + score_3_x686;
      res_4_sum <= res_4_sum + score_4_x686;
      res_5_sum <= res_5_sum + score_5_x686;
      res_6_sum <= res_6_sum + score_6_x686;
      res_7_sum <= res_7_sum + score_7_x686;
      res_8_sum <= res_8_sum + score_8_x686;
      res_9_sum <= res_9_sum + score_9_x686;
   end
   else if(res_done_x687) begin
      res_0_sum <= res_0_sum + score_0_x687;
      res_1_sum <= res_1_sum + score_1_x687;
      res_2_sum <= res_2_sum + score_2_x687;
      res_3_sum <= res_3_sum + score_3_x687;
      res_4_sum <= res_4_sum + score_4_x687;
      res_5_sum <= res_5_sum + score_5_x687;
      res_6_sum <= res_6_sum + score_6_x687;
      res_7_sum <= res_7_sum + score_7_x687;
      res_8_sum <= res_8_sum + score_8_x687;
      res_9_sum <= res_9_sum + score_9_x687;
   end
   else if(res_done_x688) begin
      res_0_sum <= res_0_sum + score_0_x688;
      res_1_sum <= res_1_sum + score_1_x688;
      res_2_sum <= res_2_sum + score_2_x688;
      res_3_sum <= res_3_sum + score_3_x688;
      res_4_sum <= res_4_sum + score_4_x688;
      res_5_sum <= res_5_sum + score_5_x688;
      res_6_sum <= res_6_sum + score_6_x688;
      res_7_sum <= res_7_sum + score_7_x688;
      res_8_sum <= res_8_sum + score_8_x688;
      res_9_sum <= res_9_sum + score_9_x688;
   end
   else if(res_done_x689) begin
      res_0_sum <= res_0_sum + score_0_x689;
      res_1_sum <= res_1_sum + score_1_x689;
      res_2_sum <= res_2_sum + score_2_x689;
      res_3_sum <= res_3_sum + score_3_x689;
      res_4_sum <= res_4_sum + score_4_x689;
      res_5_sum <= res_5_sum + score_5_x689;
      res_6_sum <= res_6_sum + score_6_x689;
      res_7_sum <= res_7_sum + score_7_x689;
      res_8_sum <= res_8_sum + score_8_x689;
      res_9_sum <= res_9_sum + score_9_x689;
   end
   else if(res_done_x690) begin
      res_0_sum <= res_0_sum + score_0_x690;
      res_1_sum <= res_1_sum + score_1_x690;
      res_2_sum <= res_2_sum + score_2_x690;
      res_3_sum <= res_3_sum + score_3_x690;
      res_4_sum <= res_4_sum + score_4_x690;
      res_5_sum <= res_5_sum + score_5_x690;
      res_6_sum <= res_6_sum + score_6_x690;
      res_7_sum <= res_7_sum + score_7_x690;
      res_8_sum <= res_8_sum + score_8_x690;
      res_9_sum <= res_9_sum + score_9_x690;
   end
   else if(res_done_x691) begin
      res_0_sum <= res_0_sum + score_0_x691;
      res_1_sum <= res_1_sum + score_1_x691;
      res_2_sum <= res_2_sum + score_2_x691;
      res_3_sum <= res_3_sum + score_3_x691;
      res_4_sum <= res_4_sum + score_4_x691;
      res_5_sum <= res_5_sum + score_5_x691;
      res_6_sum <= res_6_sum + score_6_x691;
      res_7_sum <= res_7_sum + score_7_x691;
      res_8_sum <= res_8_sum + score_8_x691;
      res_9_sum <= res_9_sum + score_9_x691;
   end
   else if(res_done_x692) begin
      res_0_sum <= res_0_sum + score_0_x692;
      res_1_sum <= res_1_sum + score_1_x692;
      res_2_sum <= res_2_sum + score_2_x692;
      res_3_sum <= res_3_sum + score_3_x692;
      res_4_sum <= res_4_sum + score_4_x692;
      res_5_sum <= res_5_sum + score_5_x692;
      res_6_sum <= res_6_sum + score_6_x692;
      res_7_sum <= res_7_sum + score_7_x692;
      res_8_sum <= res_8_sum + score_8_x692;
      res_9_sum <= res_9_sum + score_9_x692;
   end
   else if(res_done_x693) begin
      res_0_sum <= res_0_sum + score_0_x693;
      res_1_sum <= res_1_sum + score_1_x693;
      res_2_sum <= res_2_sum + score_2_x693;
      res_3_sum <= res_3_sum + score_3_x693;
      res_4_sum <= res_4_sum + score_4_x693;
      res_5_sum <= res_5_sum + score_5_x693;
      res_6_sum <= res_6_sum + score_6_x693;
      res_7_sum <= res_7_sum + score_7_x693;
      res_8_sum <= res_8_sum + score_8_x693;
      res_9_sum <= res_9_sum + score_9_x693;
   end
   else if(res_done_x694) begin
      res_0_sum <= res_0_sum + score_0_x694;
      res_1_sum <= res_1_sum + score_1_x694;
      res_2_sum <= res_2_sum + score_2_x694;
      res_3_sum <= res_3_sum + score_3_x694;
      res_4_sum <= res_4_sum + score_4_x694;
      res_5_sum <= res_5_sum + score_5_x694;
      res_6_sum <= res_6_sum + score_6_x694;
      res_7_sum <= res_7_sum + score_7_x694;
      res_8_sum <= res_8_sum + score_8_x694;
      res_9_sum <= res_9_sum + score_9_x694;
   end
   else if(res_done_x695) begin
      res_0_sum <= res_0_sum + score_0_x695;
      res_1_sum <= res_1_sum + score_1_x695;
      res_2_sum <= res_2_sum + score_2_x695;
      res_3_sum <= res_3_sum + score_3_x695;
      res_4_sum <= res_4_sum + score_4_x695;
      res_5_sum <= res_5_sum + score_5_x695;
      res_6_sum <= res_6_sum + score_6_x695;
      res_7_sum <= res_7_sum + score_7_x695;
      res_8_sum <= res_8_sum + score_8_x695;
      res_9_sum <= res_9_sum + score_9_x695;
   end
   else if(res_done_x696) begin
      res_0_sum <= res_0_sum + score_0_x696;
      res_1_sum <= res_1_sum + score_1_x696;
      res_2_sum <= res_2_sum + score_2_x696;
      res_3_sum <= res_3_sum + score_3_x696;
      res_4_sum <= res_4_sum + score_4_x696;
      res_5_sum <= res_5_sum + score_5_x696;
      res_6_sum <= res_6_sum + score_6_x696;
      res_7_sum <= res_7_sum + score_7_x696;
      res_8_sum <= res_8_sum + score_8_x696;
      res_9_sum <= res_9_sum + score_9_x696;
   end
   else if(res_done_x697) begin
      res_0_sum <= res_0_sum + score_0_x697;
      res_1_sum <= res_1_sum + score_1_x697;
      res_2_sum <= res_2_sum + score_2_x697;
      res_3_sum <= res_3_sum + score_3_x697;
      res_4_sum <= res_4_sum + score_4_x697;
      res_5_sum <= res_5_sum + score_5_x697;
      res_6_sum <= res_6_sum + score_6_x697;
      res_7_sum <= res_7_sum + score_7_x697;
      res_8_sum <= res_8_sum + score_8_x697;
      res_9_sum <= res_9_sum + score_9_x697;
   end
   else if(res_done_x698) begin
      res_0_sum <= res_0_sum + score_0_x698;
      res_1_sum <= res_1_sum + score_1_x698;
      res_2_sum <= res_2_sum + score_2_x698;
      res_3_sum <= res_3_sum + score_3_x698;
      res_4_sum <= res_4_sum + score_4_x698;
      res_5_sum <= res_5_sum + score_5_x698;
      res_6_sum <= res_6_sum + score_6_x698;
      res_7_sum <= res_7_sum + score_7_x698;
      res_8_sum <= res_8_sum + score_8_x698;
      res_9_sum <= res_9_sum + score_9_x698;
   end
   else if(res_done_x699) begin
      res_0_sum <= res_0_sum + score_0_x699;
      res_1_sum <= res_1_sum + score_1_x699;
      res_2_sum <= res_2_sum + score_2_x699;
      res_3_sum <= res_3_sum + score_3_x699;
      res_4_sum <= res_4_sum + score_4_x699;
      res_5_sum <= res_5_sum + score_5_x699;
      res_6_sum <= res_6_sum + score_6_x699;
      res_7_sum <= res_7_sum + score_7_x699;
      res_8_sum <= res_8_sum + score_8_x699;
      res_9_sum <= res_9_sum + score_9_x699;
   end
   else if(res_done_x700) begin
      res_0_sum <= res_0_sum + score_0_x700;
      res_1_sum <= res_1_sum + score_1_x700;
      res_2_sum <= res_2_sum + score_2_x700;
      res_3_sum <= res_3_sum + score_3_x700;
      res_4_sum <= res_4_sum + score_4_x700;
      res_5_sum <= res_5_sum + score_5_x700;
      res_6_sum <= res_6_sum + score_6_x700;
      res_7_sum <= res_7_sum + score_7_x700;
      res_8_sum <= res_8_sum + score_8_x700;
      res_9_sum <= res_9_sum + score_9_x700;
   end
   else if(res_done_x701) begin
      res_0_sum <= res_0_sum + score_0_x701;
      res_1_sum <= res_1_sum + score_1_x701;
      res_2_sum <= res_2_sum + score_2_x701;
      res_3_sum <= res_3_sum + score_3_x701;
      res_4_sum <= res_4_sum + score_4_x701;
      res_5_sum <= res_5_sum + score_5_x701;
      res_6_sum <= res_6_sum + score_6_x701;
      res_7_sum <= res_7_sum + score_7_x701;
      res_8_sum <= res_8_sum + score_8_x701;
      res_9_sum <= res_9_sum + score_9_x701;
   end
   else if(res_done_x702) begin
      res_0_sum <= res_0_sum + score_0_x702;
      res_1_sum <= res_1_sum + score_1_x702;
      res_2_sum <= res_2_sum + score_2_x702;
      res_3_sum <= res_3_sum + score_3_x702;
      res_4_sum <= res_4_sum + score_4_x702;
      res_5_sum <= res_5_sum + score_5_x702;
      res_6_sum <= res_6_sum + score_6_x702;
      res_7_sum <= res_7_sum + score_7_x702;
      res_8_sum <= res_8_sum + score_8_x702;
      res_9_sum <= res_9_sum + score_9_x702;
   end
   else if(res_done_x703) begin
      res_0_sum <= res_0_sum + score_0_x703;
      res_1_sum <= res_1_sum + score_1_x703;
      res_2_sum <= res_2_sum + score_2_x703;
      res_3_sum <= res_3_sum + score_3_x703;
      res_4_sum <= res_4_sum + score_4_x703;
      res_5_sum <= res_5_sum + score_5_x703;
      res_6_sum <= res_6_sum + score_6_x703;
      res_7_sum <= res_7_sum + score_7_x703;
      res_8_sum <= res_8_sum + score_8_x703;
      res_9_sum <= res_9_sum + score_9_x703;
   end
   else if(res_done_x704) begin
      res_0_sum <= res_0_sum + score_0_x704;
      res_1_sum <= res_1_sum + score_1_x704;
      res_2_sum <= res_2_sum + score_2_x704;
      res_3_sum <= res_3_sum + score_3_x704;
      res_4_sum <= res_4_sum + score_4_x704;
      res_5_sum <= res_5_sum + score_5_x704;
      res_6_sum <= res_6_sum + score_6_x704;
      res_7_sum <= res_7_sum + score_7_x704;
      res_8_sum <= res_8_sum + score_8_x704;
      res_9_sum <= res_9_sum + score_9_x704;
   end
   else if(res_done_x705) begin
      res_0_sum <= res_0_sum + score_0_x705;
      res_1_sum <= res_1_sum + score_1_x705;
      res_2_sum <= res_2_sum + score_2_x705;
      res_3_sum <= res_3_sum + score_3_x705;
      res_4_sum <= res_4_sum + score_4_x705;
      res_5_sum <= res_5_sum + score_5_x705;
      res_6_sum <= res_6_sum + score_6_x705;
      res_7_sum <= res_7_sum + score_7_x705;
      res_8_sum <= res_8_sum + score_8_x705;
      res_9_sum <= res_9_sum + score_9_x705;
   end
   else if(res_done_x706) begin
      res_0_sum <= res_0_sum + score_0_x706;
      res_1_sum <= res_1_sum + score_1_x706;
      res_2_sum <= res_2_sum + score_2_x706;
      res_3_sum <= res_3_sum + score_3_x706;
      res_4_sum <= res_4_sum + score_4_x706;
      res_5_sum <= res_5_sum + score_5_x706;
      res_6_sum <= res_6_sum + score_6_x706;
      res_7_sum <= res_7_sum + score_7_x706;
      res_8_sum <= res_8_sum + score_8_x706;
      res_9_sum <= res_9_sum + score_9_x706;
   end
   else if(res_done_x707) begin
      res_0_sum <= res_0_sum + score_0_x707;
      res_1_sum <= res_1_sum + score_1_x707;
      res_2_sum <= res_2_sum + score_2_x707;
      res_3_sum <= res_3_sum + score_3_x707;
      res_4_sum <= res_4_sum + score_4_x707;
      res_5_sum <= res_5_sum + score_5_x707;
      res_6_sum <= res_6_sum + score_6_x707;
      res_7_sum <= res_7_sum + score_7_x707;
      res_8_sum <= res_8_sum + score_8_x707;
      res_9_sum <= res_9_sum + score_9_x707;
   end
   else if(res_done_x708) begin
      res_0_sum <= res_0_sum + score_0_x708;
      res_1_sum <= res_1_sum + score_1_x708;
      res_2_sum <= res_2_sum + score_2_x708;
      res_3_sum <= res_3_sum + score_3_x708;
      res_4_sum <= res_4_sum + score_4_x708;
      res_5_sum <= res_5_sum + score_5_x708;
      res_6_sum <= res_6_sum + score_6_x708;
      res_7_sum <= res_7_sum + score_7_x708;
      res_8_sum <= res_8_sum + score_8_x708;
      res_9_sum <= res_9_sum + score_9_x708;
   end
   else if(res_done_x709) begin
      res_0_sum <= res_0_sum + score_0_x709;
      res_1_sum <= res_1_sum + score_1_x709;
      res_2_sum <= res_2_sum + score_2_x709;
      res_3_sum <= res_3_sum + score_3_x709;
      res_4_sum <= res_4_sum + score_4_x709;
      res_5_sum <= res_5_sum + score_5_x709;
      res_6_sum <= res_6_sum + score_6_x709;
      res_7_sum <= res_7_sum + score_7_x709;
      res_8_sum <= res_8_sum + score_8_x709;
      res_9_sum <= res_9_sum + score_9_x709;
   end
   else if(res_done_x710) begin
      res_0_sum <= res_0_sum + score_0_x710;
      res_1_sum <= res_1_sum + score_1_x710;
      res_2_sum <= res_2_sum + score_2_x710;
      res_3_sum <= res_3_sum + score_3_x710;
      res_4_sum <= res_4_sum + score_4_x710;
      res_5_sum <= res_5_sum + score_5_x710;
      res_6_sum <= res_6_sum + score_6_x710;
      res_7_sum <= res_7_sum + score_7_x710;
      res_8_sum <= res_8_sum + score_8_x710;
      res_9_sum <= res_9_sum + score_9_x710;
   end
   else if(res_done_x711) begin
      res_0_sum <= res_0_sum + score_0_x711;
      res_1_sum <= res_1_sum + score_1_x711;
      res_2_sum <= res_2_sum + score_2_x711;
      res_3_sum <= res_3_sum + score_3_x711;
      res_4_sum <= res_4_sum + score_4_x711;
      res_5_sum <= res_5_sum + score_5_x711;
      res_6_sum <= res_6_sum + score_6_x711;
      res_7_sum <= res_7_sum + score_7_x711;
      res_8_sum <= res_8_sum + score_8_x711;
      res_9_sum <= res_9_sum + score_9_x711;
   end
   else if(res_done_x712) begin
      res_0_sum <= res_0_sum + score_0_x712;
      res_1_sum <= res_1_sum + score_1_x712;
      res_2_sum <= res_2_sum + score_2_x712;
      res_3_sum <= res_3_sum + score_3_x712;
      res_4_sum <= res_4_sum + score_4_x712;
      res_5_sum <= res_5_sum + score_5_x712;
      res_6_sum <= res_6_sum + score_6_x712;
      res_7_sum <= res_7_sum + score_7_x712;
      res_8_sum <= res_8_sum + score_8_x712;
      res_9_sum <= res_9_sum + score_9_x712;
   end
   else if(res_done_x713) begin
      res_0_sum <= res_0_sum + score_0_x713;
      res_1_sum <= res_1_sum + score_1_x713;
      res_2_sum <= res_2_sum + score_2_x713;
      res_3_sum <= res_3_sum + score_3_x713;
      res_4_sum <= res_4_sum + score_4_x713;
      res_5_sum <= res_5_sum + score_5_x713;
      res_6_sum <= res_6_sum + score_6_x713;
      res_7_sum <= res_7_sum + score_7_x713;
      res_8_sum <= res_8_sum + score_8_x713;
      res_9_sum <= res_9_sum + score_9_x713;
   end
   else if(res_done_x714) begin
      res_0_sum <= res_0_sum + score_0_x714;
      res_1_sum <= res_1_sum + score_1_x714;
      res_2_sum <= res_2_sum + score_2_x714;
      res_3_sum <= res_3_sum + score_3_x714;
      res_4_sum <= res_4_sum + score_4_x714;
      res_5_sum <= res_5_sum + score_5_x714;
      res_6_sum <= res_6_sum + score_6_x714;
      res_7_sum <= res_7_sum + score_7_x714;
      res_8_sum <= res_8_sum + score_8_x714;
      res_9_sum <= res_9_sum + score_9_x714;
   end
   else if(res_done_x715) begin
      res_0_sum <= res_0_sum + score_0_x715;
      res_1_sum <= res_1_sum + score_1_x715;
      res_2_sum <= res_2_sum + score_2_x715;
      res_3_sum <= res_3_sum + score_3_x715;
      res_4_sum <= res_4_sum + score_4_x715;
      res_5_sum <= res_5_sum + score_5_x715;
      res_6_sum <= res_6_sum + score_6_x715;
      res_7_sum <= res_7_sum + score_7_x715;
      res_8_sum <= res_8_sum + score_8_x715;
      res_9_sum <= res_9_sum + score_9_x715;
   end
   else if(res_done_x716) begin
      res_0_sum <= res_0_sum + score_0_x716;
      res_1_sum <= res_1_sum + score_1_x716;
      res_2_sum <= res_2_sum + score_2_x716;
      res_3_sum <= res_3_sum + score_3_x716;
      res_4_sum <= res_4_sum + score_4_x716;
      res_5_sum <= res_5_sum + score_5_x716;
      res_6_sum <= res_6_sum + score_6_x716;
      res_7_sum <= res_7_sum + score_7_x716;
      res_8_sum <= res_8_sum + score_8_x716;
      res_9_sum <= res_9_sum + score_9_x716;
   end
   else if(res_done_x717) begin
      res_0_sum <= res_0_sum + score_0_x717;
      res_1_sum <= res_1_sum + score_1_x717;
      res_2_sum <= res_2_sum + score_2_x717;
      res_3_sum <= res_3_sum + score_3_x717;
      res_4_sum <= res_4_sum + score_4_x717;
      res_5_sum <= res_5_sum + score_5_x717;
      res_6_sum <= res_6_sum + score_6_x717;
      res_7_sum <= res_7_sum + score_7_x717;
      res_8_sum <= res_8_sum + score_8_x717;
      res_9_sum <= res_9_sum + score_9_x717;
   end
   else if(res_done_x718) begin
      res_0_sum <= res_0_sum + score_0_x718;
      res_1_sum <= res_1_sum + score_1_x718;
      res_2_sum <= res_2_sum + score_2_x718;
      res_3_sum <= res_3_sum + score_3_x718;
      res_4_sum <= res_4_sum + score_4_x718;
      res_5_sum <= res_5_sum + score_5_x718;
      res_6_sum <= res_6_sum + score_6_x718;
      res_7_sum <= res_7_sum + score_7_x718;
      res_8_sum <= res_8_sum + score_8_x718;
      res_9_sum <= res_9_sum + score_9_x718;
   end
   else if(res_done_x719) begin
      res_0_sum <= res_0_sum + score_0_x719;
      res_1_sum <= res_1_sum + score_1_x719;
      res_2_sum <= res_2_sum + score_2_x719;
      res_3_sum <= res_3_sum + score_3_x719;
      res_4_sum <= res_4_sum + score_4_x719;
      res_5_sum <= res_5_sum + score_5_x719;
      res_6_sum <= res_6_sum + score_6_x719;
      res_7_sum <= res_7_sum + score_7_x719;
      res_8_sum <= res_8_sum + score_8_x719;
      res_9_sum <= res_9_sum + score_9_x719;
   end
   else if(res_done_x720) begin
      res_0_sum <= res_0_sum + score_0_x720;
      res_1_sum <= res_1_sum + score_1_x720;
      res_2_sum <= res_2_sum + score_2_x720;
      res_3_sum <= res_3_sum + score_3_x720;
      res_4_sum <= res_4_sum + score_4_x720;
      res_5_sum <= res_5_sum + score_5_x720;
      res_6_sum <= res_6_sum + score_6_x720;
      res_7_sum <= res_7_sum + score_7_x720;
      res_8_sum <= res_8_sum + score_8_x720;
      res_9_sum <= res_9_sum + score_9_x720;
   end
   else if(res_done_x721) begin
      res_0_sum <= res_0_sum + score_0_x721;
      res_1_sum <= res_1_sum + score_1_x721;
      res_2_sum <= res_2_sum + score_2_x721;
      res_3_sum <= res_3_sum + score_3_x721;
      res_4_sum <= res_4_sum + score_4_x721;
      res_5_sum <= res_5_sum + score_5_x721;
      res_6_sum <= res_6_sum + score_6_x721;
      res_7_sum <= res_7_sum + score_7_x721;
      res_8_sum <= res_8_sum + score_8_x721;
      res_9_sum <= res_9_sum + score_9_x721;
   end
   else if(res_done_x722) begin
      res_0_sum <= res_0_sum + score_0_x722;
      res_1_sum <= res_1_sum + score_1_x722;
      res_2_sum <= res_2_sum + score_2_x722;
      res_3_sum <= res_3_sum + score_3_x722;
      res_4_sum <= res_4_sum + score_4_x722;
      res_5_sum <= res_5_sum + score_5_x722;
      res_6_sum <= res_6_sum + score_6_x722;
      res_7_sum <= res_7_sum + score_7_x722;
      res_8_sum <= res_8_sum + score_8_x722;
      res_9_sum <= res_9_sum + score_9_x722;
   end
   else if(res_done_x723) begin
      res_0_sum <= res_0_sum + score_0_x723;
      res_1_sum <= res_1_sum + score_1_x723;
      res_2_sum <= res_2_sum + score_2_x723;
      res_3_sum <= res_3_sum + score_3_x723;
      res_4_sum <= res_4_sum + score_4_x723;
      res_5_sum <= res_5_sum + score_5_x723;
      res_6_sum <= res_6_sum + score_6_x723;
      res_7_sum <= res_7_sum + score_7_x723;
      res_8_sum <= res_8_sum + score_8_x723;
      res_9_sum <= res_9_sum + score_9_x723;
   end
   else if(res_done_x724) begin
      res_0_sum <= res_0_sum + score_0_x724;
      res_1_sum <= res_1_sum + score_1_x724;
      res_2_sum <= res_2_sum + score_2_x724;
      res_3_sum <= res_3_sum + score_3_x724;
      res_4_sum <= res_4_sum + score_4_x724;
      res_5_sum <= res_5_sum + score_5_x724;
      res_6_sum <= res_6_sum + score_6_x724;
      res_7_sum <= res_7_sum + score_7_x724;
      res_8_sum <= res_8_sum + score_8_x724;
      res_9_sum <= res_9_sum + score_9_x724;
   end
   else if(res_done_x725) begin
      res_0_sum <= res_0_sum + score_0_x725;
      res_1_sum <= res_1_sum + score_1_x725;
      res_2_sum <= res_2_sum + score_2_x725;
      res_3_sum <= res_3_sum + score_3_x725;
      res_4_sum <= res_4_sum + score_4_x725;
      res_5_sum <= res_5_sum + score_5_x725;
      res_6_sum <= res_6_sum + score_6_x725;
      res_7_sum <= res_7_sum + score_7_x725;
      res_8_sum <= res_8_sum + score_8_x725;
      res_9_sum <= res_9_sum + score_9_x725;
   end
   else if(res_done_x726) begin
      res_0_sum <= res_0_sum + score_0_x726;
      res_1_sum <= res_1_sum + score_1_x726;
      res_2_sum <= res_2_sum + score_2_x726;
      res_3_sum <= res_3_sum + score_3_x726;
      res_4_sum <= res_4_sum + score_4_x726;
      res_5_sum <= res_5_sum + score_5_x726;
      res_6_sum <= res_6_sum + score_6_x726;
      res_7_sum <= res_7_sum + score_7_x726;
      res_8_sum <= res_8_sum + score_8_x726;
      res_9_sum <= res_9_sum + score_9_x726;
   end
   else if(res_done_x727) begin
      res_0_sum <= res_0_sum + score_0_x727;
      res_1_sum <= res_1_sum + score_1_x727;
      res_2_sum <= res_2_sum + score_2_x727;
      res_3_sum <= res_3_sum + score_3_x727;
      res_4_sum <= res_4_sum + score_4_x727;
      res_5_sum <= res_5_sum + score_5_x727;
      res_6_sum <= res_6_sum + score_6_x727;
      res_7_sum <= res_7_sum + score_7_x727;
      res_8_sum <= res_8_sum + score_8_x727;
      res_9_sum <= res_9_sum + score_9_x727;
   end
   else if(res_done_x728) begin
      res_0_sum <= res_0_sum + score_0_x728;
      res_1_sum <= res_1_sum + score_1_x728;
      res_2_sum <= res_2_sum + score_2_x728;
      res_3_sum <= res_3_sum + score_3_x728;
      res_4_sum <= res_4_sum + score_4_x728;
      res_5_sum <= res_5_sum + score_5_x728;
      res_6_sum <= res_6_sum + score_6_x728;
      res_7_sum <= res_7_sum + score_7_x728;
      res_8_sum <= res_8_sum + score_8_x728;
      res_9_sum <= res_9_sum + score_9_x728;
   end
   else if(res_done_x729) begin
      res_0_sum <= res_0_sum + score_0_x729;
      res_1_sum <= res_1_sum + score_1_x729;
      res_2_sum <= res_2_sum + score_2_x729;
      res_3_sum <= res_3_sum + score_3_x729;
      res_4_sum <= res_4_sum + score_4_x729;
      res_5_sum <= res_5_sum + score_5_x729;
      res_6_sum <= res_6_sum + score_6_x729;
      res_7_sum <= res_7_sum + score_7_x729;
      res_8_sum <= res_8_sum + score_8_x729;
      res_9_sum <= res_9_sum + score_9_x729;
   end
   else if(res_done_x730) begin
      res_0_sum <= res_0_sum + score_0_x730;
      res_1_sum <= res_1_sum + score_1_x730;
      res_2_sum <= res_2_sum + score_2_x730;
      res_3_sum <= res_3_sum + score_3_x730;
      res_4_sum <= res_4_sum + score_4_x730;
      res_5_sum <= res_5_sum + score_5_x730;
      res_6_sum <= res_6_sum + score_6_x730;
      res_7_sum <= res_7_sum + score_7_x730;
      res_8_sum <= res_8_sum + score_8_x730;
      res_9_sum <= res_9_sum + score_9_x730;
   end
   else if(res_done_x731) begin
      res_0_sum <= res_0_sum + score_0_x731;
      res_1_sum <= res_1_sum + score_1_x731;
      res_2_sum <= res_2_sum + score_2_x731;
      res_3_sum <= res_3_sum + score_3_x731;
      res_4_sum <= res_4_sum + score_4_x731;
      res_5_sum <= res_5_sum + score_5_x731;
      res_6_sum <= res_6_sum + score_6_x731;
      res_7_sum <= res_7_sum + score_7_x731;
      res_8_sum <= res_8_sum + score_8_x731;
      res_9_sum <= res_9_sum + score_9_x731;
   end
   else if(res_done_x732) begin
      res_0_sum <= res_0_sum + score_0_x732;
      res_1_sum <= res_1_sum + score_1_x732;
      res_2_sum <= res_2_sum + score_2_x732;
      res_3_sum <= res_3_sum + score_3_x732;
      res_4_sum <= res_4_sum + score_4_x732;
      res_5_sum <= res_5_sum + score_5_x732;
      res_6_sum <= res_6_sum + score_6_x732;
      res_7_sum <= res_7_sum + score_7_x732;
      res_8_sum <= res_8_sum + score_8_x732;
      res_9_sum <= res_9_sum + score_9_x732;
   end
   else if(res_done_x733) begin
      res_0_sum <= res_0_sum + score_0_x733;
      res_1_sum <= res_1_sum + score_1_x733;
      res_2_sum <= res_2_sum + score_2_x733;
      res_3_sum <= res_3_sum + score_3_x733;
      res_4_sum <= res_4_sum + score_4_x733;
      res_5_sum <= res_5_sum + score_5_x733;
      res_6_sum <= res_6_sum + score_6_x733;
      res_7_sum <= res_7_sum + score_7_x733;
      res_8_sum <= res_8_sum + score_8_x733;
      res_9_sum <= res_9_sum + score_9_x733;
   end
   else if(res_done_x734) begin
      res_0_sum <= res_0_sum + score_0_x734;
      res_1_sum <= res_1_sum + score_1_x734;
      res_2_sum <= res_2_sum + score_2_x734;
      res_3_sum <= res_3_sum + score_3_x734;
      res_4_sum <= res_4_sum + score_4_x734;
      res_5_sum <= res_5_sum + score_5_x734;
      res_6_sum <= res_6_sum + score_6_x734;
      res_7_sum <= res_7_sum + score_7_x734;
      res_8_sum <= res_8_sum + score_8_x734;
      res_9_sum <= res_9_sum + score_9_x734;
   end
   else if(res_done_x735) begin
      res_0_sum <= res_0_sum + score_0_x735;
      res_1_sum <= res_1_sum + score_1_x735;
      res_2_sum <= res_2_sum + score_2_x735;
      res_3_sum <= res_3_sum + score_3_x735;
      res_4_sum <= res_4_sum + score_4_x735;
      res_5_sum <= res_5_sum + score_5_x735;
      res_6_sum <= res_6_sum + score_6_x735;
      res_7_sum <= res_7_sum + score_7_x735;
      res_8_sum <= res_8_sum + score_8_x735;
      res_9_sum <= res_9_sum + score_9_x735;
   end
   else if(res_done_x736) begin
      res_0_sum <= res_0_sum + score_0_x736;
      res_1_sum <= res_1_sum + score_1_x736;
      res_2_sum <= res_2_sum + score_2_x736;
      res_3_sum <= res_3_sum + score_3_x736;
      res_4_sum <= res_4_sum + score_4_x736;
      res_5_sum <= res_5_sum + score_5_x736;
      res_6_sum <= res_6_sum + score_6_x736;
      res_7_sum <= res_7_sum + score_7_x736;
      res_8_sum <= res_8_sum + score_8_x736;
      res_9_sum <= res_9_sum + score_9_x736;
   end
   else if(res_done_x737) begin
      res_0_sum <= res_0_sum + score_0_x737;
      res_1_sum <= res_1_sum + score_1_x737;
      res_2_sum <= res_2_sum + score_2_x737;
      res_3_sum <= res_3_sum + score_3_x737;
      res_4_sum <= res_4_sum + score_4_x737;
      res_5_sum <= res_5_sum + score_5_x737;
      res_6_sum <= res_6_sum + score_6_x737;
      res_7_sum <= res_7_sum + score_7_x737;
      res_8_sum <= res_8_sum + score_8_x737;
      res_9_sum <= res_9_sum + score_9_x737;
   end
   else if(res_done_x738) begin
      res_0_sum <= res_0_sum + score_0_x738;
      res_1_sum <= res_1_sum + score_1_x738;
      res_2_sum <= res_2_sum + score_2_x738;
      res_3_sum <= res_3_sum + score_3_x738;
      res_4_sum <= res_4_sum + score_4_x738;
      res_5_sum <= res_5_sum + score_5_x738;
      res_6_sum <= res_6_sum + score_6_x738;
      res_7_sum <= res_7_sum + score_7_x738;
      res_8_sum <= res_8_sum + score_8_x738;
      res_9_sum <= res_9_sum + score_9_x738;
   end
   else if(res_done_x739) begin
      res_0_sum <= res_0_sum + score_0_x739;
      res_1_sum <= res_1_sum + score_1_x739;
      res_2_sum <= res_2_sum + score_2_x739;
      res_3_sum <= res_3_sum + score_3_x739;
      res_4_sum <= res_4_sum + score_4_x739;
      res_5_sum <= res_5_sum + score_5_x739;
      res_6_sum <= res_6_sum + score_6_x739;
      res_7_sum <= res_7_sum + score_7_x739;
      res_8_sum <= res_8_sum + score_8_x739;
      res_9_sum <= res_9_sum + score_9_x739;
   end
   else if(res_done_x740) begin
      res_0_sum <= res_0_sum + score_0_x740;
      res_1_sum <= res_1_sum + score_1_x740;
      res_2_sum <= res_2_sum + score_2_x740;
      res_3_sum <= res_3_sum + score_3_x740;
      res_4_sum <= res_4_sum + score_4_x740;
      res_5_sum <= res_5_sum + score_5_x740;
      res_6_sum <= res_6_sum + score_6_x740;
      res_7_sum <= res_7_sum + score_7_x740;
      res_8_sum <= res_8_sum + score_8_x740;
      res_9_sum <= res_9_sum + score_9_x740;
   end
   else if(res_done_x741) begin
      res_0_sum <= res_0_sum + score_0_x741;
      res_1_sum <= res_1_sum + score_1_x741;
      res_2_sum <= res_2_sum + score_2_x741;
      res_3_sum <= res_3_sum + score_3_x741;
      res_4_sum <= res_4_sum + score_4_x741;
      res_5_sum <= res_5_sum + score_5_x741;
      res_6_sum <= res_6_sum + score_6_x741;
      res_7_sum <= res_7_sum + score_7_x741;
      res_8_sum <= res_8_sum + score_8_x741;
      res_9_sum <= res_9_sum + score_9_x741;
   end
   else if(res_done_x742) begin
      res_0_sum <= res_0_sum + score_0_x742;
      res_1_sum <= res_1_sum + score_1_x742;
      res_2_sum <= res_2_sum + score_2_x742;
      res_3_sum <= res_3_sum + score_3_x742;
      res_4_sum <= res_4_sum + score_4_x742;
      res_5_sum <= res_5_sum + score_5_x742;
      res_6_sum <= res_6_sum + score_6_x742;
      res_7_sum <= res_7_sum + score_7_x742;
      res_8_sum <= res_8_sum + score_8_x742;
      res_9_sum <= res_9_sum + score_9_x742;
   end
   else if(res_done_x743) begin
      res_0_sum <= res_0_sum + score_0_x743;
      res_1_sum <= res_1_sum + score_1_x743;
      res_2_sum <= res_2_sum + score_2_x743;
      res_3_sum <= res_3_sum + score_3_x743;
      res_4_sum <= res_4_sum + score_4_x743;
      res_5_sum <= res_5_sum + score_5_x743;
      res_6_sum <= res_6_sum + score_6_x743;
      res_7_sum <= res_7_sum + score_7_x743;
      res_8_sum <= res_8_sum + score_8_x743;
      res_9_sum <= res_9_sum + score_9_x743;
   end
   else if(res_done_x744) begin
      res_0_sum <= res_0_sum + score_0_x744;
      res_1_sum <= res_1_sum + score_1_x744;
      res_2_sum <= res_2_sum + score_2_x744;
      res_3_sum <= res_3_sum + score_3_x744;
      res_4_sum <= res_4_sum + score_4_x744;
      res_5_sum <= res_5_sum + score_5_x744;
      res_6_sum <= res_6_sum + score_6_x744;
      res_7_sum <= res_7_sum + score_7_x744;
      res_8_sum <= res_8_sum + score_8_x744;
      res_9_sum <= res_9_sum + score_9_x744;
   end
   else if(res_done_x745) begin
      res_0_sum <= res_0_sum + score_0_x745;
      res_1_sum <= res_1_sum + score_1_x745;
      res_2_sum <= res_2_sum + score_2_x745;
      res_3_sum <= res_3_sum + score_3_x745;
      res_4_sum <= res_4_sum + score_4_x745;
      res_5_sum <= res_5_sum + score_5_x745;
      res_6_sum <= res_6_sum + score_6_x745;
      res_7_sum <= res_7_sum + score_7_x745;
      res_8_sum <= res_8_sum + score_8_x745;
      res_9_sum <= res_9_sum + score_9_x745;
   end
   else if(res_done_x746) begin
      res_0_sum <= res_0_sum + score_0_x746;
      res_1_sum <= res_1_sum + score_1_x746;
      res_2_sum <= res_2_sum + score_2_x746;
      res_3_sum <= res_3_sum + score_3_x746;
      res_4_sum <= res_4_sum + score_4_x746;
      res_5_sum <= res_5_sum + score_5_x746;
      res_6_sum <= res_6_sum + score_6_x746;
      res_7_sum <= res_7_sum + score_7_x746;
      res_8_sum <= res_8_sum + score_8_x746;
      res_9_sum <= res_9_sum + score_9_x746;
   end
   else if(res_done_x747) begin
      res_0_sum <= res_0_sum + score_0_x747;
      res_1_sum <= res_1_sum + score_1_x747;
      res_2_sum <= res_2_sum + score_2_x747;
      res_3_sum <= res_3_sum + score_3_x747;
      res_4_sum <= res_4_sum + score_4_x747;
      res_5_sum <= res_5_sum + score_5_x747;
      res_6_sum <= res_6_sum + score_6_x747;
      res_7_sum <= res_7_sum + score_7_x747;
      res_8_sum <= res_8_sum + score_8_x747;
      res_9_sum <= res_9_sum + score_9_x747;
   end
   else if(res_done_x748) begin
      res_0_sum <= res_0_sum + score_0_x748;
      res_1_sum <= res_1_sum + score_1_x748;
      res_2_sum <= res_2_sum + score_2_x748;
      res_3_sum <= res_3_sum + score_3_x748;
      res_4_sum <= res_4_sum + score_4_x748;
      res_5_sum <= res_5_sum + score_5_x748;
      res_6_sum <= res_6_sum + score_6_x748;
      res_7_sum <= res_7_sum + score_7_x748;
      res_8_sum <= res_8_sum + score_8_x748;
      res_9_sum <= res_9_sum + score_9_x748;
   end
   else if(res_done_x749) begin
      res_0_sum <= res_0_sum + score_0_x749;
      res_1_sum <= res_1_sum + score_1_x749;
      res_2_sum <= res_2_sum + score_2_x749;
      res_3_sum <= res_3_sum + score_3_x749;
      res_4_sum <= res_4_sum + score_4_x749;
      res_5_sum <= res_5_sum + score_5_x749;
      res_6_sum <= res_6_sum + score_6_x749;
      res_7_sum <= res_7_sum + score_7_x749;
      res_8_sum <= res_8_sum + score_8_x749;
      res_9_sum <= res_9_sum + score_9_x749;
   end
   else if(res_done_x750) begin
      res_0_sum <= res_0_sum + score_0_x750;
      res_1_sum <= res_1_sum + score_1_x750;
      res_2_sum <= res_2_sum + score_2_x750;
      res_3_sum <= res_3_sum + score_3_x750;
      res_4_sum <= res_4_sum + score_4_x750;
      res_5_sum <= res_5_sum + score_5_x750;
      res_6_sum <= res_6_sum + score_6_x750;
      res_7_sum <= res_7_sum + score_7_x750;
      res_8_sum <= res_8_sum + score_8_x750;
      res_9_sum <= res_9_sum + score_9_x750;
   end
   else if(res_done_x751) begin
      res_0_sum <= res_0_sum + score_0_x751;
      res_1_sum <= res_1_sum + score_1_x751;
      res_2_sum <= res_2_sum + score_2_x751;
      res_3_sum <= res_3_sum + score_3_x751;
      res_4_sum <= res_4_sum + score_4_x751;
      res_5_sum <= res_5_sum + score_5_x751;
      res_6_sum <= res_6_sum + score_6_x751;
      res_7_sum <= res_7_sum + score_7_x751;
      res_8_sum <= res_8_sum + score_8_x751;
      res_9_sum <= res_9_sum + score_9_x751;
   end
   else if(res_done_x752) begin
      res_0_sum <= res_0_sum + score_0_x752;
      res_1_sum <= res_1_sum + score_1_x752;
      res_2_sum <= res_2_sum + score_2_x752;
      res_3_sum <= res_3_sum + score_3_x752;
      res_4_sum <= res_4_sum + score_4_x752;
      res_5_sum <= res_5_sum + score_5_x752;
      res_6_sum <= res_6_sum + score_6_x752;
      res_7_sum <= res_7_sum + score_7_x752;
      res_8_sum <= res_8_sum + score_8_x752;
      res_9_sum <= res_9_sum + score_9_x752;
   end
   else if(res_done_x753) begin
      res_0_sum <= res_0_sum + score_0_x753;
      res_1_sum <= res_1_sum + score_1_x753;
      res_2_sum <= res_2_sum + score_2_x753;
      res_3_sum <= res_3_sum + score_3_x753;
      res_4_sum <= res_4_sum + score_4_x753;
      res_5_sum <= res_5_sum + score_5_x753;
      res_6_sum <= res_6_sum + score_6_x753;
      res_7_sum <= res_7_sum + score_7_x753;
      res_8_sum <= res_8_sum + score_8_x753;
      res_9_sum <= res_9_sum + score_9_x753;
   end
   else if(res_done_x754) begin
      res_0_sum <= res_0_sum + score_0_x754;
      res_1_sum <= res_1_sum + score_1_x754;
      res_2_sum <= res_2_sum + score_2_x754;
      res_3_sum <= res_3_sum + score_3_x754;
      res_4_sum <= res_4_sum + score_4_x754;
      res_5_sum <= res_5_sum + score_5_x754;
      res_6_sum <= res_6_sum + score_6_x754;
      res_7_sum <= res_7_sum + score_7_x754;
      res_8_sum <= res_8_sum + score_8_x754;
      res_9_sum <= res_9_sum + score_9_x754;
   end
   else if(res_done_x755) begin
      res_0_sum <= res_0_sum + score_0_x755;
      res_1_sum <= res_1_sum + score_1_x755;
      res_2_sum <= res_2_sum + score_2_x755;
      res_3_sum <= res_3_sum + score_3_x755;
      res_4_sum <= res_4_sum + score_4_x755;
      res_5_sum <= res_5_sum + score_5_x755;
      res_6_sum <= res_6_sum + score_6_x755;
      res_7_sum <= res_7_sum + score_7_x755;
      res_8_sum <= res_8_sum + score_8_x755;
      res_9_sum <= res_9_sum + score_9_x755;
   end
   else if(res_done_x756) begin
      res_0_sum <= res_0_sum + score_0_x756;
      res_1_sum <= res_1_sum + score_1_x756;
      res_2_sum <= res_2_sum + score_2_x756;
      res_3_sum <= res_3_sum + score_3_x756;
      res_4_sum <= res_4_sum + score_4_x756;
      res_5_sum <= res_5_sum + score_5_x756;
      res_6_sum <= res_6_sum + score_6_x756;
      res_7_sum <= res_7_sum + score_7_x756;
      res_8_sum <= res_8_sum + score_8_x756;
      res_9_sum <= res_9_sum + score_9_x756;
   end
   else if(res_done_x757) begin
      res_0_sum <= res_0_sum + score_0_x757;
      res_1_sum <= res_1_sum + score_1_x757;
      res_2_sum <= res_2_sum + score_2_x757;
      res_3_sum <= res_3_sum + score_3_x757;
      res_4_sum <= res_4_sum + score_4_x757;
      res_5_sum <= res_5_sum + score_5_x757;
      res_6_sum <= res_6_sum + score_6_x757;
      res_7_sum <= res_7_sum + score_7_x757;
      res_8_sum <= res_8_sum + score_8_x757;
      res_9_sum <= res_9_sum + score_9_x757;
   end
   else if(res_done_x758) begin
      res_0_sum <= res_0_sum + score_0_x758;
      res_1_sum <= res_1_sum + score_1_x758;
      res_2_sum <= res_2_sum + score_2_x758;
      res_3_sum <= res_3_sum + score_3_x758;
      res_4_sum <= res_4_sum + score_4_x758;
      res_5_sum <= res_5_sum + score_5_x758;
      res_6_sum <= res_6_sum + score_6_x758;
      res_7_sum <= res_7_sum + score_7_x758;
      res_8_sum <= res_8_sum + score_8_x758;
      res_9_sum <= res_9_sum + score_9_x758;
   end
   else if(res_done_x759) begin
      res_0_sum <= res_0_sum + score_0_x759;
      res_1_sum <= res_1_sum + score_1_x759;
      res_2_sum <= res_2_sum + score_2_x759;
      res_3_sum <= res_3_sum + score_3_x759;
      res_4_sum <= res_4_sum + score_4_x759;
      res_5_sum <= res_5_sum + score_5_x759;
      res_6_sum <= res_6_sum + score_6_x759;
      res_7_sum <= res_7_sum + score_7_x759;
      res_8_sum <= res_8_sum + score_8_x759;
      res_9_sum <= res_9_sum + score_9_x759;
   end
   else if(res_done_x760) begin
      res_0_sum <= res_0_sum + score_0_x760;
      res_1_sum <= res_1_sum + score_1_x760;
      res_2_sum <= res_2_sum + score_2_x760;
      res_3_sum <= res_3_sum + score_3_x760;
      res_4_sum <= res_4_sum + score_4_x760;
      res_5_sum <= res_5_sum + score_5_x760;
      res_6_sum <= res_6_sum + score_6_x760;
      res_7_sum <= res_7_sum + score_7_x760;
      res_8_sum <= res_8_sum + score_8_x760;
      res_9_sum <= res_9_sum + score_9_x760;
   end
   else if(res_done_x761) begin
      res_0_sum <= res_0_sum + score_0_x761;
      res_1_sum <= res_1_sum + score_1_x761;
      res_2_sum <= res_2_sum + score_2_x761;
      res_3_sum <= res_3_sum + score_3_x761;
      res_4_sum <= res_4_sum + score_4_x761;
      res_5_sum <= res_5_sum + score_5_x761;
      res_6_sum <= res_6_sum + score_6_x761;
      res_7_sum <= res_7_sum + score_7_x761;
      res_8_sum <= res_8_sum + score_8_x761;
      res_9_sum <= res_9_sum + score_9_x761;
   end
   else if(res_done_x762) begin
      res_0_sum <= res_0_sum + score_0_x762;
      res_1_sum <= res_1_sum + score_1_x762;
      res_2_sum <= res_2_sum + score_2_x762;
      res_3_sum <= res_3_sum + score_3_x762;
      res_4_sum <= res_4_sum + score_4_x762;
      res_5_sum <= res_5_sum + score_5_x762;
      res_6_sum <= res_6_sum + score_6_x762;
      res_7_sum <= res_7_sum + score_7_x762;
      res_8_sum <= res_8_sum + score_8_x762;
      res_9_sum <= res_9_sum + score_9_x762;
   end
   else if(res_done_x763) begin
      res_0_sum <= res_0_sum + score_0_x763;
      res_1_sum <= res_1_sum + score_1_x763;
      res_2_sum <= res_2_sum + score_2_x763;
      res_3_sum <= res_3_sum + score_3_x763;
      res_4_sum <= res_4_sum + score_4_x763;
      res_5_sum <= res_5_sum + score_5_x763;
      res_6_sum <= res_6_sum + score_6_x763;
      res_7_sum <= res_7_sum + score_7_x763;
      res_8_sum <= res_8_sum + score_8_x763;
      res_9_sum <= res_9_sum + score_9_x763;
   end
   else if(res_done_x764) begin
      res_0_sum <= res_0_sum + score_0_x764;
      res_1_sum <= res_1_sum + score_1_x764;
      res_2_sum <= res_2_sum + score_2_x764;
      res_3_sum <= res_3_sum + score_3_x764;
      res_4_sum <= res_4_sum + score_4_x764;
      res_5_sum <= res_5_sum + score_5_x764;
      res_6_sum <= res_6_sum + score_6_x764;
      res_7_sum <= res_7_sum + score_7_x764;
      res_8_sum <= res_8_sum + score_8_x764;
      res_9_sum <= res_9_sum + score_9_x764;
   end
   else if(res_done_x765) begin
      res_0_sum <= res_0_sum + score_0_x765;
      res_1_sum <= res_1_sum + score_1_x765;
      res_2_sum <= res_2_sum + score_2_x765;
      res_3_sum <= res_3_sum + score_3_x765;
      res_4_sum <= res_4_sum + score_4_x765;
      res_5_sum <= res_5_sum + score_5_x765;
      res_6_sum <= res_6_sum + score_6_x765;
      res_7_sum <= res_7_sum + score_7_x765;
      res_8_sum <= res_8_sum + score_8_x765;
      res_9_sum <= res_9_sum + score_9_x765;
   end
   else if(res_done_x766) begin
      res_0_sum <= res_0_sum + score_0_x766;
      res_1_sum <= res_1_sum + score_1_x766;
      res_2_sum <= res_2_sum + score_2_x766;
      res_3_sum <= res_3_sum + score_3_x766;
      res_4_sum <= res_4_sum + score_4_x766;
      res_5_sum <= res_5_sum + score_5_x766;
      res_6_sum <= res_6_sum + score_6_x766;
      res_7_sum <= res_7_sum + score_7_x766;
      res_8_sum <= res_8_sum + score_8_x766;
      res_9_sum <= res_9_sum + score_9_x766;
   end
   else if(res_done_x767) begin
      res_0_sum <= res_0_sum + score_0_x767;
      res_1_sum <= res_1_sum + score_1_x767;
      res_2_sum <= res_2_sum + score_2_x767;
      res_3_sum <= res_3_sum + score_3_x767;
      res_4_sum <= res_4_sum + score_4_x767;
      res_5_sum <= res_5_sum + score_5_x767;
      res_6_sum <= res_6_sum + score_6_x767;
      res_7_sum <= res_7_sum + score_7_x767;
      res_8_sum <= res_8_sum + score_8_x767;
      res_9_sum <= res_9_sum + score_9_x767;
   end
   else if(res_done_x768) begin
      res_0_sum <= res_0_sum + score_0_x768;
      res_1_sum <= res_1_sum + score_1_x768;
      res_2_sum <= res_2_sum + score_2_x768;
      res_3_sum <= res_3_sum + score_3_x768;
      res_4_sum <= res_4_sum + score_4_x768;
      res_5_sum <= res_5_sum + score_5_x768;
      res_6_sum <= res_6_sum + score_6_x768;
      res_7_sum <= res_7_sum + score_7_x768;
      res_8_sum <= res_8_sum + score_8_x768;
      res_9_sum <= res_9_sum + score_9_x768;
   end
   else if(res_done_x769) begin
      res_0_sum <= res_0_sum + score_0_x769;
      res_1_sum <= res_1_sum + score_1_x769;
      res_2_sum <= res_2_sum + score_2_x769;
      res_3_sum <= res_3_sum + score_3_x769;
      res_4_sum <= res_4_sum + score_4_x769;
      res_5_sum <= res_5_sum + score_5_x769;
      res_6_sum <= res_6_sum + score_6_x769;
      res_7_sum <= res_7_sum + score_7_x769;
      res_8_sum <= res_8_sum + score_8_x769;
      res_9_sum <= res_9_sum + score_9_x769;
   end
   else if(res_done_x770) begin
      res_0_sum <= res_0_sum + score_0_x770;
      res_1_sum <= res_1_sum + score_1_x770;
      res_2_sum <= res_2_sum + score_2_x770;
      res_3_sum <= res_3_sum + score_3_x770;
      res_4_sum <= res_4_sum + score_4_x770;
      res_5_sum <= res_5_sum + score_5_x770;
      res_6_sum <= res_6_sum + score_6_x770;
      res_7_sum <= res_7_sum + score_7_x770;
      res_8_sum <= res_8_sum + score_8_x770;
      res_9_sum <= res_9_sum + score_9_x770;
   end
   else if(res_done_x771) begin
      res_0_sum <= res_0_sum + score_0_x771;
      res_1_sum <= res_1_sum + score_1_x771;
      res_2_sum <= res_2_sum + score_2_x771;
      res_3_sum <= res_3_sum + score_3_x771;
      res_4_sum <= res_4_sum + score_4_x771;
      res_5_sum <= res_5_sum + score_5_x771;
      res_6_sum <= res_6_sum + score_6_x771;
      res_7_sum <= res_7_sum + score_7_x771;
      res_8_sum <= res_8_sum + score_8_x771;
      res_9_sum <= res_9_sum + score_9_x771;
   end
   else if(res_done_x772) begin
      res_0_sum <= res_0_sum + score_0_x772;
      res_1_sum <= res_1_sum + score_1_x772;
      res_2_sum <= res_2_sum + score_2_x772;
      res_3_sum <= res_3_sum + score_3_x772;
      res_4_sum <= res_4_sum + score_4_x772;
      res_5_sum <= res_5_sum + score_5_x772;
      res_6_sum <= res_6_sum + score_6_x772;
      res_7_sum <= res_7_sum + score_7_x772;
      res_8_sum <= res_8_sum + score_8_x772;
      res_9_sum <= res_9_sum + score_9_x772;
   end
   else if(res_done_x773) begin
      res_0_sum <= res_0_sum + score_0_x773;
      res_1_sum <= res_1_sum + score_1_x773;
      res_2_sum <= res_2_sum + score_2_x773;
      res_3_sum <= res_3_sum + score_3_x773;
      res_4_sum <= res_4_sum + score_4_x773;
      res_5_sum <= res_5_sum + score_5_x773;
      res_6_sum <= res_6_sum + score_6_x773;
      res_7_sum <= res_7_sum + score_7_x773;
      res_8_sum <= res_8_sum + score_8_x773;
      res_9_sum <= res_9_sum + score_9_x773;
   end
   else if(res_done_x774) begin
      res_0_sum <= res_0_sum + score_0_x774;
      res_1_sum <= res_1_sum + score_1_x774;
      res_2_sum <= res_2_sum + score_2_x774;
      res_3_sum <= res_3_sum + score_3_x774;
      res_4_sum <= res_4_sum + score_4_x774;
      res_5_sum <= res_5_sum + score_5_x774;
      res_6_sum <= res_6_sum + score_6_x774;
      res_7_sum <= res_7_sum + score_7_x774;
      res_8_sum <= res_8_sum + score_8_x774;
      res_9_sum <= res_9_sum + score_9_x774;
   end
   else if(res_done_x775) begin
      res_0_sum <= res_0_sum + score_0_x775;
      res_1_sum <= res_1_sum + score_1_x775;
      res_2_sum <= res_2_sum + score_2_x775;
      res_3_sum <= res_3_sum + score_3_x775;
      res_4_sum <= res_4_sum + score_4_x775;
      res_5_sum <= res_5_sum + score_5_x775;
      res_6_sum <= res_6_sum + score_6_x775;
      res_7_sum <= res_7_sum + score_7_x775;
      res_8_sum <= res_8_sum + score_8_x775;
      res_9_sum <= res_9_sum + score_9_x775;
   end
   else if(res_done_x776) begin
      res_0_sum <= res_0_sum + score_0_x776;
      res_1_sum <= res_1_sum + score_1_x776;
      res_2_sum <= res_2_sum + score_2_x776;
      res_3_sum <= res_3_sum + score_3_x776;
      res_4_sum <= res_4_sum + score_4_x776;
      res_5_sum <= res_5_sum + score_5_x776;
      res_6_sum <= res_6_sum + score_6_x776;
      res_7_sum <= res_7_sum + score_7_x776;
      res_8_sum <= res_8_sum + score_8_x776;
      res_9_sum <= res_9_sum + score_9_x776;
   end
   else if(res_done_x777) begin
      res_0_sum <= res_0_sum + score_0_x777;
      res_1_sum <= res_1_sum + score_1_x777;
      res_2_sum <= res_2_sum + score_2_x777;
      res_3_sum <= res_3_sum + score_3_x777;
      res_4_sum <= res_4_sum + score_4_x777;
      res_5_sum <= res_5_sum + score_5_x777;
      res_6_sum <= res_6_sum + score_6_x777;
      res_7_sum <= res_7_sum + score_7_x777;
      res_8_sum <= res_8_sum + score_8_x777;
      res_9_sum <= res_9_sum + score_9_x777;
   end
   else if(res_done_x778) begin
      res_0_sum <= res_0_sum + score_0_x778;
      res_1_sum <= res_1_sum + score_1_x778;
      res_2_sum <= res_2_sum + score_2_x778;
      res_3_sum <= res_3_sum + score_3_x778;
      res_4_sum <= res_4_sum + score_4_x778;
      res_5_sum <= res_5_sum + score_5_x778;
      res_6_sum <= res_6_sum + score_6_x778;
      res_7_sum <= res_7_sum + score_7_x778;
      res_8_sum <= res_8_sum + score_8_x778;
      res_9_sum <= res_9_sum + score_9_x778;
   end
   else if(res_done_x779) begin
      res_0_sum <= res_0_sum + score_0_x779;
      res_1_sum <= res_1_sum + score_1_x779;
      res_2_sum <= res_2_sum + score_2_x779;
      res_3_sum <= res_3_sum + score_3_x779;
      res_4_sum <= res_4_sum + score_4_x779;
      res_5_sum <= res_5_sum + score_5_x779;
      res_6_sum <= res_6_sum + score_6_x779;
      res_7_sum <= res_7_sum + score_7_x779;
      res_8_sum <= res_8_sum + score_8_x779;
      res_9_sum <= res_9_sum + score_9_x779;
   end
   else if(res_done_x780) begin
      res_0_sum <= res_0_sum + score_0_x780;
      res_1_sum <= res_1_sum + score_1_x780;
      res_2_sum <= res_2_sum + score_2_x780;
      res_3_sum <= res_3_sum + score_3_x780;
      res_4_sum <= res_4_sum + score_4_x780;
      res_5_sum <= res_5_sum + score_5_x780;
      res_6_sum <= res_6_sum + score_6_x780;
      res_7_sum <= res_7_sum + score_7_x780;
      res_8_sum <= res_8_sum + score_8_x780;
      res_9_sum <= res_9_sum + score_9_x780;
   end
   else if(res_done_x781) begin
      res_0_sum <= res_0_sum + score_0_x781;
      res_1_sum <= res_1_sum + score_1_x781;
      res_2_sum <= res_2_sum + score_2_x781;
      res_3_sum <= res_3_sum + score_3_x781;
      res_4_sum <= res_4_sum + score_4_x781;
      res_5_sum <= res_5_sum + score_5_x781;
      res_6_sum <= res_6_sum + score_6_x781;
      res_7_sum <= res_7_sum + score_7_x781;
      res_8_sum <= res_8_sum + score_8_x781;
      res_9_sum <= res_9_sum + score_9_x781;
   end
   else if(res_done_x782) begin
      res_0_sum <= res_0_sum + score_0_x782;
      res_1_sum <= res_1_sum + score_1_x782;
      res_2_sum <= res_2_sum + score_2_x782;
      res_3_sum <= res_3_sum + score_3_x782;
      res_4_sum <= res_4_sum + score_4_x782;
      res_5_sum <= res_5_sum + score_5_x782;
      res_6_sum <= res_6_sum + score_6_x782;
      res_7_sum <= res_7_sum + score_7_x782;
      res_8_sum <= res_8_sum + score_8_x782;
      res_9_sum <= res_9_sum + score_9_x782;
   end
   else if(res_done_x783) begin
      res_0_sum <= res_0_sum + score_0_x783;
      res_1_sum <= res_1_sum + score_1_x783;
      res_2_sum <= res_2_sum + score_2_x783;
      res_3_sum <= res_3_sum + score_3_x783;
      res_4_sum <= res_4_sum + score_4_x783;
      res_5_sum <= res_5_sum + score_5_x783;
      res_6_sum <= res_6_sum + score_6_x783;
      res_7_sum <= res_7_sum + score_7_x783;
      res_8_sum <= res_8_sum + score_8_x783;
      res_9_sum <= res_9_sum + score_9_x783;
   end
   else if(res_done_x784) begin
      res_0_sum <= res_0_sum + score_0_x784;
      res_1_sum <= res_1_sum + score_1_x784;
      res_2_sum <= res_2_sum + score_2_x784;
      res_3_sum <= res_3_sum + score_3_x784;
      res_4_sum <= res_4_sum + score_4_x784;
      res_5_sum <= res_5_sum + score_5_x784;
      res_6_sum <= res_6_sum + score_6_x784;
      res_7_sum <= res_7_sum + score_7_x784;
      res_8_sum <= res_8_sum + score_8_x784;
      res_9_sum <= res_9_sum + score_9_x784;
   end
   else if(done_all_res[1]) begin	
        res_0_sum <= res_0_sum + B_0;
        res_1_sum <= res_1_sum + B_1;
        res_2_sum <= res_2_sum + B_2;
        res_3_sum <= res_3_sum + B_3;
        res_4_sum <= res_4_sum + B_4;
        res_5_sum <= res_5_sum + B_5;
        res_6_sum <= res_6_sum + B_6;
        res_7_sum <= res_7_sum + B_7;
        res_8_sum <= res_8_sum + B_8;
        res_9_sum <= res_9_sum + B_9;
    end 
    else begin
    	res_0_sum <= res_0_sum;
        res_1_sum <= res_1_sum;
        res_2_sum <= res_2_sum;
        res_3_sum <= res_3_sum;
        res_4_sum <= res_4_sum;
        res_5_sum <= res_5_sum;
        res_6_sum <= res_6_sum;
        res_7_sum <= res_7_sum;
        res_8_sum <= res_8_sum;
        res_9_sum <= res_9_sum;



    end 

end







//****************************    W 输入    *******************************

localparam signed [DEBIT:0]  W_0_x1 =  23'd962;
localparam signed [DEBIT:0]  W_0_x2 =  23'd969;
localparam signed [DEBIT:0]  W_0_x3 =  23'd972;
localparam signed [DEBIT:0]  W_0_x4 =  23'd975;
localparam signed [DEBIT:0]  W_0_x5 =  23'd973;
localparam signed [DEBIT:0]  W_0_x6 =  23'd969;
localparam signed [DEBIT:0]  W_0_x7 =  23'd973;
localparam signed [DEBIT:0]  W_0_x8 =  23'd969;
localparam signed [DEBIT:0]  W_0_x9 =  23'd964;
localparam signed [DEBIT:0]  W_0_x10 =  23'd973;
localparam signed [DEBIT:0]  W_0_x11 =  23'd973;
localparam signed [DEBIT:0]  W_0_x12 =  23'd961;
localparam signed [DEBIT:0]  W_0_x13 =  23'd967;
localparam signed [DEBIT:0]  W_0_x14 =  23'd966;
localparam signed [DEBIT:0]  W_0_x15 =  23'd966;
localparam signed [DEBIT:0]  W_0_x16 =  23'd959;
localparam signed [DEBIT:0]  W_0_x17 =  23'd968;
localparam signed [DEBIT:0]  W_0_x18 =  23'd975;
localparam signed [DEBIT:0]  W_0_x19 =  23'd968;
localparam signed [DEBIT:0]  W_0_x20 =  23'd961;
localparam signed [DEBIT:0]  W_0_x21 =  23'd969;
localparam signed [DEBIT:0]  W_0_x22 =  23'd960;
localparam signed [DEBIT:0]  W_0_x23 =  23'd977;
localparam signed [DEBIT:0]  W_0_x24 =  23'd966;
localparam signed [DEBIT:0]  W_0_x25 =  23'd968;
localparam signed [DEBIT:0]  W_0_x26 =  23'd970;
localparam signed [DEBIT:0]  W_0_x27 =  23'd958;
localparam signed [DEBIT:0]  W_0_x28 =  23'd958;
localparam signed [DEBIT:0]  W_0_x29 =  23'd971;
localparam signed [DEBIT:0]  W_0_x30 =  23'd962;
localparam signed [DEBIT:0]  W_0_x31 =  23'd959;
localparam signed [DEBIT:0]  W_0_x32 =  23'd961;
localparam signed [DEBIT:0]  W_0_x33 =  23'd963;
localparam signed [DEBIT:0]  W_0_x34 =  23'd967;
localparam signed [DEBIT:0]  W_0_x35 =  23'd973;
localparam signed [DEBIT:0]  W_0_x36 =  23'd975;
localparam signed [DEBIT:0]  W_0_x37 =  23'd968;
localparam signed [DEBIT:0]  W_0_x38 =  23'd953;
localparam signed [DEBIT:0]  W_0_x39 =  23'd960;
localparam signed [DEBIT:0]  W_0_x40 =  23'd968;
localparam signed [DEBIT:0]  W_0_x41 =  23'd963;
localparam signed [DEBIT:0]  W_0_x42 =  23'd960;
localparam signed [DEBIT:0]  W_0_x43 =  23'd953;
localparam signed [DEBIT:0]  W_0_x44 =  23'd955;
localparam signed [DEBIT:0]  W_0_x45 =  23'd951;
localparam signed [DEBIT:0]  W_0_x46 =  23'd950;
localparam signed [DEBIT:0]  W_0_x47 =  23'd969;
localparam signed [DEBIT:0]  W_0_x48 =  23'd964;
localparam signed [DEBIT:0]  W_0_x49 =  23'd960;
localparam signed [DEBIT:0]  W_0_x50 =  23'd967;
localparam signed [DEBIT:0]  W_0_x51 =  23'd973;
localparam signed [DEBIT:0]  W_0_x52 =  23'd964;
localparam signed [DEBIT:0]  W_0_x53 =  23'd965;
localparam signed [DEBIT:0]  W_0_x54 =  23'd960;
localparam signed [DEBIT:0]  W_0_x55 =  23'd970;
localparam signed [DEBIT:0]  W_0_x56 =  23'd964;
localparam signed [DEBIT:0]  W_0_x57 =  23'd975;
localparam signed [DEBIT:0]  W_0_x58 =  23'd968;
localparam signed [DEBIT:0]  W_0_x59 =  23'd971;
localparam signed [DEBIT:0]  W_0_x60 =  23'd965;
localparam signed [DEBIT:0]  W_0_x61 =  23'd971;
localparam signed [DEBIT:0]  W_0_x62 =  23'd967;
localparam signed [DEBIT:0]  W_0_x63 =  23'd962;
localparam signed [DEBIT:0]  W_0_x64 =  23'd937;
localparam signed [DEBIT:0]  W_0_x65 =  23'd894;
localparam signed [DEBIT:0]  W_0_x66 =  23'd815;
localparam signed [DEBIT:0]  W_0_x67 =  23'd829;
localparam signed [DEBIT:0]  W_0_x68 =  23'd836;
localparam signed [DEBIT:0]  W_0_x69 =  23'd780;
localparam signed [DEBIT:0]  W_0_x70 =  23'd757;
localparam signed [DEBIT:0]  W_0_x71 =  23'd704;
localparam signed [DEBIT:0]  W_0_x72 =  23'd693;
localparam signed [DEBIT:0]  W_0_x73 =  23'd687;
localparam signed [DEBIT:0]  W_0_x74 =  23'd755;
localparam signed [DEBIT:0]  W_0_x75 =  23'd791;
localparam signed [DEBIT:0]  W_0_x76 =  23'd785;
localparam signed [DEBIT:0]  W_0_x77 =  23'd844;
localparam signed [DEBIT:0]  W_0_x78 =  23'd894;
localparam signed [DEBIT:0]  W_0_x79 =  23'd914;
localparam signed [DEBIT:0]  W_0_x80 =  23'd943;
localparam signed [DEBIT:0]  W_0_x81 =  23'd966;
localparam signed [DEBIT:0]  W_0_x82 =  23'd953;
localparam signed [DEBIT:0]  W_0_x83 =  23'd962;
localparam signed [DEBIT:0]  W_0_x84 =  23'd966;
localparam signed [DEBIT:0]  W_0_x85 =  23'd968;
localparam signed [DEBIT:0]  W_0_x86 =  23'd974;
localparam signed [DEBIT:0]  W_0_x87 =  23'd960;
localparam signed [DEBIT:0]  W_0_x88 =  23'd962;
localparam signed [DEBIT:0]  W_0_x89 =  23'd978;
localparam signed [DEBIT:0]  W_0_x90 =  23'd942;
localparam signed [DEBIT:0]  W_0_x91 =  23'd898;
localparam signed [DEBIT:0]  W_0_x92 =  23'd815;
localparam signed [DEBIT:0]  W_0_x93 =  23'd652;
localparam signed [DEBIT:0]  W_0_x94 =  23'd525;
localparam signed [DEBIT:0]  W_0_x95 =  23'd440;
localparam signed [DEBIT:0]  W_0_x96 =  23'd366;
localparam signed [DEBIT:0]  W_0_x97 =  23'd294;
localparam signed [DEBIT:0]  W_0_x98 =  23'd261;
localparam signed [DEBIT:0]  W_0_x99 =  23'd170;
localparam signed [DEBIT:0]  W_0_x100 =  23'd151;
localparam signed [DEBIT:0]  W_0_x101 =  23'd171;
localparam signed [DEBIT:0]  W_0_x102 =  23'd257;
localparam signed [DEBIT:0]  W_0_x103 =  23'd305;
localparam signed [DEBIT:0]  W_0_x104 =  23'd366;
localparam signed [DEBIT:0]  W_0_x105 =  23'd484;
localparam signed [DEBIT:0]  W_0_x106 =  23'd616;
localparam signed [DEBIT:0]  W_0_x107 =  23'd753;
localparam signed [DEBIT:0]  W_0_x108 =  23'd869;
localparam signed [DEBIT:0]  W_0_x109 =  23'd939;
localparam signed [DEBIT:0]  W_0_x110 =  23'd972;
localparam signed [DEBIT:0]  W_0_x111 =  23'd968;
localparam signed [DEBIT:0]  W_0_x112 =  23'd972;
localparam signed [DEBIT:0]  W_0_x113 =  23'd969;
localparam signed [DEBIT:0]  W_0_x114 =  23'd972;
localparam signed [DEBIT:0]  W_0_x115 =  23'd977;
localparam signed [DEBIT:0]  W_0_x116 =  23'd956;
localparam signed [DEBIT:0]  W_0_x117 =  23'd951;
localparam signed [DEBIT:0]  W_0_x118 =  23'd871;
localparam signed [DEBIT:0]  W_0_x119 =  23'd763;
localparam signed [DEBIT:0]  W_0_x120 =  23'd562;
localparam signed [DEBIT:0]  W_0_x121 =  23'd333;
localparam signed [DEBIT:0]  W_0_x122 =  23'd164;
localparam signed [DEBIT:0]  W_0_x123 =  23'd107;
localparam signed [DEBIT:0]  W_0_x124 =  23'd52;
localparam signed [DEBIT:0]  W_0_x125 =  23'd25;
localparam signed [DEBIT:0]  W_0_x126 =  23'd69;
localparam signed [DEBIT:0]  W_0_x127 =  23'd111;
localparam signed [DEBIT:0]  W_0_x128 =  23'd84;
localparam signed [DEBIT:0]  W_0_x129 =  23'd22;
localparam signed [DEBIT:0]  W_0_x130 =  23'd119;
localparam signed [DEBIT:0]  W_0_x131 =  23'd133;
localparam signed [DEBIT:0]  W_0_x132 =  23'd99;
localparam signed [DEBIT:0]  W_0_x133 =  23'd154;
localparam signed [DEBIT:0]  W_0_x134 =  23'd281;
localparam signed [DEBIT:0]  W_0_x135 =  23'd434;
localparam signed [DEBIT:0]  W_0_x136 =  23'd683;
localparam signed [DEBIT:0]  W_0_x137 =  23'd827;
localparam signed [DEBIT:0]  W_0_x138 =  23'd923;
localparam signed [DEBIT:0]  W_0_x139 =  23'd964;
localparam signed [DEBIT:0]  W_0_x140 =  23'd970;
localparam signed [DEBIT:0]  W_0_x141 =  23'd962;
localparam signed [DEBIT:0]  W_0_x142 =  23'd968;
localparam signed [DEBIT:0]  W_0_x143 =  23'd964;
localparam signed [DEBIT:0]  W_0_x144 =  23'd963;
localparam signed [DEBIT:0]  W_0_x145 =  23'd901;
localparam signed [DEBIT:0]  W_0_x146 =  23'd716;
localparam signed [DEBIT:0]  W_0_x147 =  23'd458;
localparam signed [DEBIT:0]  W_0_x148 =  23'd168;
localparam signed [DEBIT:0]  W_0_x149 = - 23'd26;
localparam signed [DEBIT:0]  W_0_x150 = - 23'd153;
localparam signed [DEBIT:0]  W_0_x151 = - 23'd124;
localparam signed [DEBIT:0]  W_0_x152 = - 23'd84;
localparam signed [DEBIT:0]  W_0_x153 =  23'd71;
localparam signed [DEBIT:0]  W_0_x154 =  23'd100;
localparam signed [DEBIT:0]  W_0_x155 =  23'd206;
localparam signed [DEBIT:0]  W_0_x156 =  23'd181;
localparam signed [DEBIT:0]  W_0_x157 =  23'd112;
localparam signed [DEBIT:0]  W_0_x158 =  23'd77;
localparam signed [DEBIT:0]  W_0_x159 =  23'd65;
localparam signed [DEBIT:0]  W_0_x160 = - 23'd2;
localparam signed [DEBIT:0]  W_0_x161 = - 23'd77;
localparam signed [DEBIT:0]  W_0_x162 = - 23'd100;
localparam signed [DEBIT:0]  W_0_x163 =  23'd130;
localparam signed [DEBIT:0]  W_0_x164 =  23'd392;
localparam signed [DEBIT:0]  W_0_x165 =  23'd604;
localparam signed [DEBIT:0]  W_0_x166 =  23'd805;
localparam signed [DEBIT:0]  W_0_x167 =  23'd937;
localparam signed [DEBIT:0]  W_0_x168 =  23'd964;
localparam signed [DEBIT:0]  W_0_x169 =  23'd973;
localparam signed [DEBIT:0]  W_0_x170 =  23'd968;
localparam signed [DEBIT:0]  W_0_x171 =  23'd967;
localparam signed [DEBIT:0]  W_0_x172 =  23'd926;
localparam signed [DEBIT:0]  W_0_x173 =  23'd778;
localparam signed [DEBIT:0]  W_0_x174 =  23'd554;
localparam signed [DEBIT:0]  W_0_x175 =  23'd278;
localparam signed [DEBIT:0]  W_0_x176 =  23'd20;
localparam signed [DEBIT:0]  W_0_x177 = - 23'd181;
localparam signed [DEBIT:0]  W_0_x178 = - 23'd271;
localparam signed [DEBIT:0]  W_0_x179 = - 23'd139;
localparam signed [DEBIT:0]  W_0_x180 =  23'd13;
localparam signed [DEBIT:0]  W_0_x181 =  23'd129;
localparam signed [DEBIT:0]  W_0_x182 =  23'd184;
localparam signed [DEBIT:0]  W_0_x183 =  23'd216;
localparam signed [DEBIT:0]  W_0_x184 =  23'd195;
localparam signed [DEBIT:0]  W_0_x185 =  23'd252;
localparam signed [DEBIT:0]  W_0_x186 =  23'd272;
localparam signed [DEBIT:0]  W_0_x187 =  23'd173;
localparam signed [DEBIT:0]  W_0_x188 =  23'd81;
localparam signed [DEBIT:0]  W_0_x189 = - 23'd164;
localparam signed [DEBIT:0]  W_0_x190 = - 23'd251;
localparam signed [DEBIT:0]  W_0_x191 = - 23'd139;
localparam signed [DEBIT:0]  W_0_x192 =  23'd153;
localparam signed [DEBIT:0]  W_0_x193 =  23'd368;
localparam signed [DEBIT:0]  W_0_x194 =  23'd628;
localparam signed [DEBIT:0]  W_0_x195 =  23'd852;
localparam signed [DEBIT:0]  W_0_x196 =  23'd943;
localparam signed [DEBIT:0]  W_0_x197 =  23'd972;
localparam signed [DEBIT:0]  W_0_x198 =  23'd960;
localparam signed [DEBIT:0]  W_0_x199 =  23'd932;
localparam signed [DEBIT:0]  W_0_x200 =  23'd847;
localparam signed [DEBIT:0]  W_0_x201 =  23'd630;
localparam signed [DEBIT:0]  W_0_x202 =  23'd362;
localparam signed [DEBIT:0]  W_0_x203 =  23'd85;
localparam signed [DEBIT:0]  W_0_x204 = - 23'd176;
localparam signed [DEBIT:0]  W_0_x205 = - 23'd230;
localparam signed [DEBIT:0]  W_0_x206 = - 23'd135;
localparam signed [DEBIT:0]  W_0_x207 =  23'd37;
localparam signed [DEBIT:0]  W_0_x208 =  23'd135;
localparam signed [DEBIT:0]  W_0_x209 =  23'd138;
localparam signed [DEBIT:0]  W_0_x210 =  23'd103;
localparam signed [DEBIT:0]  W_0_x211 =  23'd151;
localparam signed [DEBIT:0]  W_0_x212 =  23'd213;
localparam signed [DEBIT:0]  W_0_x213 =  23'd243;
localparam signed [DEBIT:0]  W_0_x214 =  23'd394;
localparam signed [DEBIT:0]  W_0_x215 =  23'd328;
localparam signed [DEBIT:0]  W_0_x216 =  23'd181;
localparam signed [DEBIT:0]  W_0_x217 = - 23'd102;
localparam signed [DEBIT:0]  W_0_x218 = - 23'd283;
localparam signed [DEBIT:0]  W_0_x219 = - 23'd245;
localparam signed [DEBIT:0]  W_0_x220 = - 23'd10;
localparam signed [DEBIT:0]  W_0_x221 =  23'd252;
localparam signed [DEBIT:0]  W_0_x222 =  23'd559;
localparam signed [DEBIT:0]  W_0_x223 =  23'd857;
localparam signed [DEBIT:0]  W_0_x224 =  23'd952;
localparam signed [DEBIT:0]  W_0_x225 =  23'd968;
localparam signed [DEBIT:0]  W_0_x226 =  23'd943;
localparam signed [DEBIT:0]  W_0_x227 =  23'd865;
localparam signed [DEBIT:0]  W_0_x228 =  23'd688;
localparam signed [DEBIT:0]  W_0_x229 =  23'd356;
localparam signed [DEBIT:0]  W_0_x230 =  23'd114;
localparam signed [DEBIT:0]  W_0_x231 = - 23'd177;
localparam signed [DEBIT:0]  W_0_x232 = - 23'd394;
localparam signed [DEBIT:0]  W_0_x233 = - 23'd367;
localparam signed [DEBIT:0]  W_0_x234 = - 23'd102;
localparam signed [DEBIT:0]  W_0_x235 =  23'd18;
localparam signed [DEBIT:0]  W_0_x236 =  23'd32;
localparam signed [DEBIT:0]  W_0_x237 = - 23'd32;
localparam signed [DEBIT:0]  W_0_x238 = - 23'd94;
localparam signed [DEBIT:0]  W_0_x239 = - 23'd56;
localparam signed [DEBIT:0]  W_0_x240 =  23'd81;
localparam signed [DEBIT:0]  W_0_x241 =  23'd214;
localparam signed [DEBIT:0]  W_0_x242 =  23'd274;
localparam signed [DEBIT:0]  W_0_x243 =  23'd125;
localparam signed [DEBIT:0]  W_0_x244 =  23'd3;
localparam signed [DEBIT:0]  W_0_x245 = - 23'd83;
localparam signed [DEBIT:0]  W_0_x246 = - 23'd231;
localparam signed [DEBIT:0]  W_0_x247 = - 23'd166;
localparam signed [DEBIT:0]  W_0_x248 =  23'd74;
localparam signed [DEBIT:0]  W_0_x249 =  23'd347;
localparam signed [DEBIT:0]  W_0_x250 =  23'd572;
localparam signed [DEBIT:0]  W_0_x251 =  23'd865;
localparam signed [DEBIT:0]  W_0_x252 =  23'd960;
localparam signed [DEBIT:0]  W_0_x253 =  23'd969;
localparam signed [DEBIT:0]  W_0_x254 =  23'd914;
localparam signed [DEBIT:0]  W_0_x255 =  23'd804;
localparam signed [DEBIT:0]  W_0_x256 =  23'd583;
localparam signed [DEBIT:0]  W_0_x257 =  23'd267;
localparam signed [DEBIT:0]  W_0_x258 = - 23'd49;
localparam signed [DEBIT:0]  W_0_x259 = - 23'd368;
localparam signed [DEBIT:0]  W_0_x260 = - 23'd473;
localparam signed [DEBIT:0]  W_0_x261 = - 23'd312;
localparam signed [DEBIT:0]  W_0_x262 = - 23'd196;
localparam signed [DEBIT:0]  W_0_x263 = - 23'd97;
localparam signed [DEBIT:0]  W_0_x264 = - 23'd115;
localparam signed [DEBIT:0]  W_0_x265 = - 23'd111;
localparam signed [DEBIT:0]  W_0_x266 = - 23'd140;
localparam signed [DEBIT:0]  W_0_x267 = - 23'd119;
localparam signed [DEBIT:0]  W_0_x268 =  23'd11;
localparam signed [DEBIT:0]  W_0_x269 =  23'd138;
localparam signed [DEBIT:0]  W_0_x270 =  23'd183;
localparam signed [DEBIT:0]  W_0_x271 =  23'd148;
localparam signed [DEBIT:0]  W_0_x272 =  23'd68;
localparam signed [DEBIT:0]  W_0_x273 =  23'd45;
localparam signed [DEBIT:0]  W_0_x274 = - 23'd111;
localparam signed [DEBIT:0]  W_0_x275 = - 23'd115;
localparam signed [DEBIT:0]  W_0_x276 =  23'd160;
localparam signed [DEBIT:0]  W_0_x277 =  23'd448;
localparam signed [DEBIT:0]  W_0_x278 =  23'd636;
localparam signed [DEBIT:0]  W_0_x279 =  23'd851;
localparam signed [DEBIT:0]  W_0_x280 =  23'd957;
localparam signed [DEBIT:0]  W_0_x281 =  23'd973;
localparam signed [DEBIT:0]  W_0_x282 =  23'd905;
localparam signed [DEBIT:0]  W_0_x283 =  23'd786;
localparam signed [DEBIT:0]  W_0_x284 =  23'd571;
localparam signed [DEBIT:0]  W_0_x285 =  23'd251;
localparam signed [DEBIT:0]  W_0_x286 = - 23'd106;
localparam signed [DEBIT:0]  W_0_x287 = - 23'd392;
localparam signed [DEBIT:0]  W_0_x288 = - 23'd333;
localparam signed [DEBIT:0]  W_0_x289 = - 23'd188;
localparam signed [DEBIT:0]  W_0_x290 = - 23'd134;
localparam signed [DEBIT:0]  W_0_x291 = - 23'd221;
localparam signed [DEBIT:0]  W_0_x292 = - 23'd159;
localparam signed [DEBIT:0]  W_0_x293 = - 23'd28;
localparam signed [DEBIT:0]  W_0_x294 = - 23'd112;
localparam signed [DEBIT:0]  W_0_x295 = - 23'd178;
localparam signed [DEBIT:0]  W_0_x296 = - 23'd109;
localparam signed [DEBIT:0]  W_0_x297 = - 23'd138;
localparam signed [DEBIT:0]  W_0_x298 =  23'd204;
localparam signed [DEBIT:0]  W_0_x299 =  23'd178;
localparam signed [DEBIT:0]  W_0_x300 =  23'd118;
localparam signed [DEBIT:0]  W_0_x301 =  23'd152;
localparam signed [DEBIT:0]  W_0_x302 =  23'd128;
localparam signed [DEBIT:0]  W_0_x303 =  23'd52;
localparam signed [DEBIT:0]  W_0_x304 =  23'd303;
localparam signed [DEBIT:0]  W_0_x305 =  23'd542;
localparam signed [DEBIT:0]  W_0_x306 =  23'd713;
localparam signed [DEBIT:0]  W_0_x307 =  23'd864;
localparam signed [DEBIT:0]  W_0_x308 =  23'd948;
localparam signed [DEBIT:0]  W_0_x309 =  23'd963;
localparam signed [DEBIT:0]  W_0_x310 =  23'd914;
localparam signed [DEBIT:0]  W_0_x311 =  23'd810;
localparam signed [DEBIT:0]  W_0_x312 =  23'd583;
localparam signed [DEBIT:0]  W_0_x313 =  23'd253;
localparam signed [DEBIT:0]  W_0_x314 = - 23'd90;
localparam signed [DEBIT:0]  W_0_x315 = - 23'd278;
localparam signed [DEBIT:0]  W_0_x316 = - 23'd146;
localparam signed [DEBIT:0]  W_0_x317 = - 23'd24;
localparam signed [DEBIT:0]  W_0_x318 = - 23'd70;
localparam signed [DEBIT:0]  W_0_x319 = - 23'd93;
localparam signed [DEBIT:0]  W_0_x320 = - 23'd16;
localparam signed [DEBIT:0]  W_0_x321 = - 23'd54;
localparam signed [DEBIT:0]  W_0_x322 = - 23'd177;
localparam signed [DEBIT:0]  W_0_x323 = - 23'd395;
localparam signed [DEBIT:0]  W_0_x324 = - 23'd405;
localparam signed [DEBIT:0]  W_0_x325 = - 23'd288;
localparam signed [DEBIT:0]  W_0_x326 =  23'd63;
localparam signed [DEBIT:0]  W_0_x327 =  23'd173;
localparam signed [DEBIT:0]  W_0_x328 =  23'd163;
localparam signed [DEBIT:0]  W_0_x329 =  23'd149;
localparam signed [DEBIT:0]  W_0_x330 =  23'd180;
localparam signed [DEBIT:0]  W_0_x331 =  23'd168;
localparam signed [DEBIT:0]  W_0_x332 =  23'd416;
localparam signed [DEBIT:0]  W_0_x333 =  23'd613;
localparam signed [DEBIT:0]  W_0_x334 =  23'd804;
localparam signed [DEBIT:0]  W_0_x335 =  23'd915;
localparam signed [DEBIT:0]  W_0_x336 =  23'd960;
localparam signed [DEBIT:0]  W_0_x337 =  23'd978;
localparam signed [DEBIT:0]  W_0_x338 =  23'd956;
localparam signed [DEBIT:0]  W_0_x339 =  23'd855;
localparam signed [DEBIT:0]  W_0_x340 =  23'd646;
localparam signed [DEBIT:0]  W_0_x341 =  23'd306;
localparam signed [DEBIT:0]  W_0_x342 =  23'd46;
localparam signed [DEBIT:0]  W_0_x343 = - 23'd88;
localparam signed [DEBIT:0]  W_0_x344 = - 23'd54;
localparam signed [DEBIT:0]  W_0_x345 =  23'd141;
localparam signed [DEBIT:0]  W_0_x346 =  23'd32;
localparam signed [DEBIT:0]  W_0_x347 =  23'd2;
localparam signed [DEBIT:0]  W_0_x348 = - 23'd48;
localparam signed [DEBIT:0]  W_0_x349 = - 23'd59;
localparam signed [DEBIT:0]  W_0_x350 = - 23'd273;
localparam signed [DEBIT:0]  W_0_x351 = - 23'd584;
localparam signed [DEBIT:0]  W_0_x352 = - 23'd676;
localparam signed [DEBIT:0]  W_0_x353 = - 23'd506;
localparam signed [DEBIT:0]  W_0_x354 = - 23'd152;
localparam signed [DEBIT:0]  W_0_x355 =  23'd11;
localparam signed [DEBIT:0]  W_0_x356 = - 23'd69;
localparam signed [DEBIT:0]  W_0_x357 = - 23'd13;
localparam signed [DEBIT:0]  W_0_x358 =  23'd171;
localparam signed [DEBIT:0]  W_0_x359 =  23'd289;
localparam signed [DEBIT:0]  W_0_x360 =  23'd477;
localparam signed [DEBIT:0]  W_0_x361 =  23'd652;
localparam signed [DEBIT:0]  W_0_x362 =  23'd861;
localparam signed [DEBIT:0]  W_0_x363 =  23'd948;
localparam signed [DEBIT:0]  W_0_x364 =  23'd966;
localparam signed [DEBIT:0]  W_0_x365 =  23'd972;
localparam signed [DEBIT:0]  W_0_x366 =  23'd972;
localparam signed [DEBIT:0]  W_0_x367 =  23'd910;
localparam signed [DEBIT:0]  W_0_x368 =  23'd724;
localparam signed [DEBIT:0]  W_0_x369 =  23'd411;
localparam signed [DEBIT:0]  W_0_x370 =  23'd261;
localparam signed [DEBIT:0]  W_0_x371 =  23'd136;
localparam signed [DEBIT:0]  W_0_x372 =  23'd87;
localparam signed [DEBIT:0]  W_0_x373 =  23'd164;
localparam signed [DEBIT:0]  W_0_x374 =  23'd152;
localparam signed [DEBIT:0]  W_0_x375 =  23'd162;
localparam signed [DEBIT:0]  W_0_x376 =  23'd51;
localparam signed [DEBIT:0]  W_0_x377 =  23'd30;
localparam signed [DEBIT:0]  W_0_x378 = - 23'd391;
localparam signed [DEBIT:0]  W_0_x379 = - 23'd647;
localparam signed [DEBIT:0]  W_0_x380 = - 23'd663;
localparam signed [DEBIT:0]  W_0_x381 = - 23'd464;
localparam signed [DEBIT:0]  W_0_x382 = - 23'd271;
localparam signed [DEBIT:0]  W_0_x383 = - 23'd244;
localparam signed [DEBIT:0]  W_0_x384 = - 23'd333;
localparam signed [DEBIT:0]  W_0_x385 = - 23'd190;
localparam signed [DEBIT:0]  W_0_x386 =  23'd104;
localparam signed [DEBIT:0]  W_0_x387 =  23'd303;
localparam signed [DEBIT:0]  W_0_x388 =  23'd446;
localparam signed [DEBIT:0]  W_0_x389 =  23'd590;
localparam signed [DEBIT:0]  W_0_x390 =  23'd857;
localparam signed [DEBIT:0]  W_0_x391 =  23'd958;
localparam signed [DEBIT:0]  W_0_x392 =  23'd961;
localparam signed [DEBIT:0]  W_0_x393 =  23'd969;
localparam signed [DEBIT:0]  W_0_x394 =  23'd972;
localparam signed [DEBIT:0]  W_0_x395 =  23'd940;
localparam signed [DEBIT:0]  W_0_x396 =  23'd782;
localparam signed [DEBIT:0]  W_0_x397 =  23'd515;
localparam signed [DEBIT:0]  W_0_x398 =  23'd409;
localparam signed [DEBIT:0]  W_0_x399 =  23'd215;
localparam signed [DEBIT:0]  W_0_x400 =  23'd214;
localparam signed [DEBIT:0]  W_0_x401 =  23'd135;
localparam signed [DEBIT:0]  W_0_x402 =  23'd204;
localparam signed [DEBIT:0]  W_0_x403 =  23'd226;
localparam signed [DEBIT:0]  W_0_x404 =  23'd116;
localparam signed [DEBIT:0]  W_0_x405 = - 23'd144;
localparam signed [DEBIT:0]  W_0_x406 = - 23'd476;
localparam signed [DEBIT:0]  W_0_x407 = - 23'd557;
localparam signed [DEBIT:0]  W_0_x408 = - 23'd551;
localparam signed [DEBIT:0]  W_0_x409 = - 23'd487;
localparam signed [DEBIT:0]  W_0_x410 = - 23'd349;
localparam signed [DEBIT:0]  W_0_x411 = - 23'd258;
localparam signed [DEBIT:0]  W_0_x412 = - 23'd273;
localparam signed [DEBIT:0]  W_0_x413 = - 23'd76;
localparam signed [DEBIT:0]  W_0_x414 =  23'd96;
localparam signed [DEBIT:0]  W_0_x415 =  23'd197;
localparam signed [DEBIT:0]  W_0_x416 =  23'd390;
localparam signed [DEBIT:0]  W_0_x417 =  23'd578;
localparam signed [DEBIT:0]  W_0_x418 =  23'd825;
localparam signed [DEBIT:0]  W_0_x419 =  23'd944;
localparam signed [DEBIT:0]  W_0_x420 =  23'd967;
localparam signed [DEBIT:0]  W_0_x421 =  23'd963;
localparam signed [DEBIT:0]  W_0_x422 =  23'd966;
localparam signed [DEBIT:0]  W_0_x423 =  23'd975;
localparam signed [DEBIT:0]  W_0_x424 =  23'd787;
localparam signed [DEBIT:0]  W_0_x425 =  23'd571;
localparam signed [DEBIT:0]  W_0_x426 =  23'd452;
localparam signed [DEBIT:0]  W_0_x427 =  23'd184;
localparam signed [DEBIT:0]  W_0_x428 =  23'd215;
localparam signed [DEBIT:0]  W_0_x429 =  23'd205;
localparam signed [DEBIT:0]  W_0_x430 =  23'd316;
localparam signed [DEBIT:0]  W_0_x431 =  23'd236;
localparam signed [DEBIT:0]  W_0_x432 = - 23'd103;
localparam signed [DEBIT:0]  W_0_x433 = - 23'd404;
localparam signed [DEBIT:0]  W_0_x434 = - 23'd633;
localparam signed [DEBIT:0]  W_0_x435 = - 23'd583;
localparam signed [DEBIT:0]  W_0_x436 = - 23'd506;
localparam signed [DEBIT:0]  W_0_x437 = - 23'd485;
localparam signed [DEBIT:0]  W_0_x438 = - 23'd322;
localparam signed [DEBIT:0]  W_0_x439 = - 23'd245;
localparam signed [DEBIT:0]  W_0_x440 = - 23'd173;
localparam signed [DEBIT:0]  W_0_x441 = - 23'd16;
localparam signed [DEBIT:0]  W_0_x442 =  23'd16;
localparam signed [DEBIT:0]  W_0_x443 =  23'd109;
localparam signed [DEBIT:0]  W_0_x444 =  23'd300;
localparam signed [DEBIT:0]  W_0_x445 =  23'd498;
localparam signed [DEBIT:0]  W_0_x446 =  23'd781;
localparam signed [DEBIT:0]  W_0_x447 =  23'd939;
localparam signed [DEBIT:0]  W_0_x448 =  23'd964;
localparam signed [DEBIT:0]  W_0_x449 =  23'd971;
localparam signed [DEBIT:0]  W_0_x450 =  23'd976;
localparam signed [DEBIT:0]  W_0_x451 =  23'd952;
localparam signed [DEBIT:0]  W_0_x452 =  23'd776;
localparam signed [DEBIT:0]  W_0_x453 =  23'd554;
localparam signed [DEBIT:0]  W_0_x454 =  23'd383;
localparam signed [DEBIT:0]  W_0_x455 =  23'd190;
localparam signed [DEBIT:0]  W_0_x456 =  23'd222;
localparam signed [DEBIT:0]  W_0_x457 =  23'd305;
localparam signed [DEBIT:0]  W_0_x458 =  23'd294;
localparam signed [DEBIT:0]  W_0_x459 =  23'd270;
localparam signed [DEBIT:0]  W_0_x460 = - 23'd232;
localparam signed [DEBIT:0]  W_0_x461 = - 23'd631;
localparam signed [DEBIT:0]  W_0_x462 = - 23'd677;
localparam signed [DEBIT:0]  W_0_x463 = - 23'd617;
localparam signed [DEBIT:0]  W_0_x464 = - 23'd517;
localparam signed [DEBIT:0]  W_0_x465 = - 23'd424;
localparam signed [DEBIT:0]  W_0_x466 = - 23'd188;
localparam signed [DEBIT:0]  W_0_x467 = - 23'd159;
localparam signed [DEBIT:0]  W_0_x468 = - 23'd89;
localparam signed [DEBIT:0]  W_0_x469 =  23'd12;
localparam signed [DEBIT:0]  W_0_x470 =  23'd63;
localparam signed [DEBIT:0]  W_0_x471 =  23'd61;
localparam signed [DEBIT:0]  W_0_x472 =  23'd159;
localparam signed [DEBIT:0]  W_0_x473 =  23'd424;
localparam signed [DEBIT:0]  W_0_x474 =  23'd759;
localparam signed [DEBIT:0]  W_0_x475 =  23'd949;
localparam signed [DEBIT:0]  W_0_x476 =  23'd961;
localparam signed [DEBIT:0]  W_0_x477 =  23'd957;
localparam signed [DEBIT:0]  W_0_x478 =  23'd962;
localparam signed [DEBIT:0]  W_0_x479 =  23'd946;
localparam signed [DEBIT:0]  W_0_x480 =  23'd759;
localparam signed [DEBIT:0]  W_0_x481 =  23'd480;
localparam signed [DEBIT:0]  W_0_x482 =  23'd331;
localparam signed [DEBIT:0]  W_0_x483 =  23'd276;
localparam signed [DEBIT:0]  W_0_x484 =  23'd265;
localparam signed [DEBIT:0]  W_0_x485 =  23'd312;
localparam signed [DEBIT:0]  W_0_x486 =  23'd428;
localparam signed [DEBIT:0]  W_0_x487 =  23'd375;
localparam signed [DEBIT:0]  W_0_x488 = - 23'd142;
localparam signed [DEBIT:0]  W_0_x489 = - 23'd482;
localparam signed [DEBIT:0]  W_0_x490 = - 23'd710;
localparam signed [DEBIT:0]  W_0_x491 = - 23'd691;
localparam signed [DEBIT:0]  W_0_x492 = - 23'd522;
localparam signed [DEBIT:0]  W_0_x493 = - 23'd243;
localparam signed [DEBIT:0]  W_0_x494 = - 23'd73;
localparam signed [DEBIT:0]  W_0_x495 = - 23'd142;
localparam signed [DEBIT:0]  W_0_x496 = - 23'd69;
localparam signed [DEBIT:0]  W_0_x497 = - 23'd123;
localparam signed [DEBIT:0]  W_0_x498 = - 23'd63;
localparam signed [DEBIT:0]  W_0_x499 = - 23'd13;
localparam signed [DEBIT:0]  W_0_x500 =  23'd58;
localparam signed [DEBIT:0]  W_0_x501 =  23'd401;
localparam signed [DEBIT:0]  W_0_x502 =  23'd775;
localparam signed [DEBIT:0]  W_0_x503 =  23'd947;
localparam signed [DEBIT:0]  W_0_x504 =  23'd964;
localparam signed [DEBIT:0]  W_0_x505 =  23'd973;
localparam signed [DEBIT:0]  W_0_x506 =  23'd959;
localparam signed [DEBIT:0]  W_0_x507 =  23'd931;
localparam signed [DEBIT:0]  W_0_x508 =  23'd692;
localparam signed [DEBIT:0]  W_0_x509 =  23'd379;
localparam signed [DEBIT:0]  W_0_x510 =  23'd203;
localparam signed [DEBIT:0]  W_0_x511 =  23'd233;
localparam signed [DEBIT:0]  W_0_x512 =  23'd326;
localparam signed [DEBIT:0]  W_0_x513 =  23'd378;
localparam signed [DEBIT:0]  W_0_x514 =  23'd390;
localparam signed [DEBIT:0]  W_0_x515 =  23'd358;
localparam signed [DEBIT:0]  W_0_x516 =  23'd124;
localparam signed [DEBIT:0]  W_0_x517 = - 23'd340;
localparam signed [DEBIT:0]  W_0_x518 = - 23'd646;
localparam signed [DEBIT:0]  W_0_x519 = - 23'd615;
localparam signed [DEBIT:0]  W_0_x520 = - 23'd418;
localparam signed [DEBIT:0]  W_0_x521 = - 23'd259;
localparam signed [DEBIT:0]  W_0_x522 = - 23'd187;
localparam signed [DEBIT:0]  W_0_x523 = - 23'd242;
localparam signed [DEBIT:0]  W_0_x524 = - 23'd156;
localparam signed [DEBIT:0]  W_0_x525 = - 23'd204;
localparam signed [DEBIT:0]  W_0_x526 = - 23'd296;
localparam signed [DEBIT:0]  W_0_x527 = - 23'd271;
localparam signed [DEBIT:0]  W_0_x528 = - 23'd69;
localparam signed [DEBIT:0]  W_0_x529 =  23'd428;
localparam signed [DEBIT:0]  W_0_x530 =  23'd814;
localparam signed [DEBIT:0]  W_0_x531 =  23'd933;
localparam signed [DEBIT:0]  W_0_x532 =  23'd965;
localparam signed [DEBIT:0]  W_0_x533 =  23'd968;
localparam signed [DEBIT:0]  W_0_x534 =  23'd958;
localparam signed [DEBIT:0]  W_0_x535 =  23'd914;
localparam signed [DEBIT:0]  W_0_x536 =  23'd591;
localparam signed [DEBIT:0]  W_0_x537 =  23'd225;
localparam signed [DEBIT:0]  W_0_x538 =  23'd99;
localparam signed [DEBIT:0]  W_0_x539 =  23'd12;
localparam signed [DEBIT:0]  W_0_x540 =  23'd151;
localparam signed [DEBIT:0]  W_0_x541 =  23'd279;
localparam signed [DEBIT:0]  W_0_x542 =  23'd301;
localparam signed [DEBIT:0]  W_0_x543 =  23'd372;
localparam signed [DEBIT:0]  W_0_x544 =  23'd280;
localparam signed [DEBIT:0]  W_0_x545 = - 23'd50;
localparam signed [DEBIT:0]  W_0_x546 = - 23'd320;
localparam signed [DEBIT:0]  W_0_x547 = - 23'd352;
localparam signed [DEBIT:0]  W_0_x548 = - 23'd345;
localparam signed [DEBIT:0]  W_0_x549 = - 23'd286;
localparam signed [DEBIT:0]  W_0_x550 = - 23'd337;
localparam signed [DEBIT:0]  W_0_x551 = - 23'd395;
localparam signed [DEBIT:0]  W_0_x552 = - 23'd376;
localparam signed [DEBIT:0]  W_0_x553 = - 23'd330;
localparam signed [DEBIT:0]  W_0_x554 = - 23'd425;
localparam signed [DEBIT:0]  W_0_x555 = - 23'd362;
localparam signed [DEBIT:0]  W_0_x556 = - 23'd1;
localparam signed [DEBIT:0]  W_0_x557 =  23'd559;
localparam signed [DEBIT:0]  W_0_x558 =  23'd823;
localparam signed [DEBIT:0]  W_0_x559 =  23'd936;
localparam signed [DEBIT:0]  W_0_x560 =  23'd958;
localparam signed [DEBIT:0]  W_0_x561 =  23'd971;
localparam signed [DEBIT:0]  W_0_x562 =  23'd957;
localparam signed [DEBIT:0]  W_0_x563 =  23'd899;
localparam signed [DEBIT:0]  W_0_x564 =  23'd582;
localparam signed [DEBIT:0]  W_0_x565 =  23'd159;
localparam signed [DEBIT:0]  W_0_x566 =  23'd38;
localparam signed [DEBIT:0]  W_0_x567 = - 23'd112;
localparam signed [DEBIT:0]  W_0_x568 = - 23'd76;
localparam signed [DEBIT:0]  W_0_x569 = - 23'd9;
localparam signed [DEBIT:0]  W_0_x570 =  23'd123;
localparam signed [DEBIT:0]  W_0_x571 =  23'd288;
localparam signed [DEBIT:0]  W_0_x572 =  23'd263;
localparam signed [DEBIT:0]  W_0_x573 =  23'd89;
localparam signed [DEBIT:0]  W_0_x574 = - 23'd110;
localparam signed [DEBIT:0]  W_0_x575 = - 23'd263;
localparam signed [DEBIT:0]  W_0_x576 = - 23'd301;
localparam signed [DEBIT:0]  W_0_x577 = - 23'd312;
localparam signed [DEBIT:0]  W_0_x578 = - 23'd286;
localparam signed [DEBIT:0]  W_0_x579 = - 23'd390;
localparam signed [DEBIT:0]  W_0_x580 = - 23'd386;
localparam signed [DEBIT:0]  W_0_x581 = - 23'd418;
localparam signed [DEBIT:0]  W_0_x582 = - 23'd481;
localparam signed [DEBIT:0]  W_0_x583 = - 23'd306;
localparam signed [DEBIT:0]  W_0_x584 =  23'd147;
localparam signed [DEBIT:0]  W_0_x585 =  23'd614;
localparam signed [DEBIT:0]  W_0_x586 =  23'd871;
localparam signed [DEBIT:0]  W_0_x587 =  23'd959;
localparam signed [DEBIT:0]  W_0_x588 =  23'd981;
localparam signed [DEBIT:0]  W_0_x589 =  23'd966;
localparam signed [DEBIT:0]  W_0_x590 =  23'd948;
localparam signed [DEBIT:0]  W_0_x591 =  23'd890;
localparam signed [DEBIT:0]  W_0_x592 =  23'd653;
localparam signed [DEBIT:0]  W_0_x593 =  23'd288;
localparam signed [DEBIT:0]  W_0_x594 =  23'd71;
localparam signed [DEBIT:0]  W_0_x595 = - 23'd133;
localparam signed [DEBIT:0]  W_0_x596 = - 23'd217;
localparam signed [DEBIT:0]  W_0_x597 = - 23'd50;
localparam signed [DEBIT:0]  W_0_x598 =  23'd61;
localparam signed [DEBIT:0]  W_0_x599 =  23'd233;
localparam signed [DEBIT:0]  W_0_x600 =  23'd293;
localparam signed [DEBIT:0]  W_0_x601 =  23'd46;
localparam signed [DEBIT:0]  W_0_x602 = - 23'd75;
localparam signed [DEBIT:0]  W_0_x603 = - 23'd141;
localparam signed [DEBIT:0]  W_0_x604 = - 23'd160;
localparam signed [DEBIT:0]  W_0_x605 = - 23'd203;
localparam signed [DEBIT:0]  W_0_x606 = - 23'd234;
localparam signed [DEBIT:0]  W_0_x607 = - 23'd236;
localparam signed [DEBIT:0]  W_0_x608 = - 23'd355;
localparam signed [DEBIT:0]  W_0_x609 = - 23'd462;
localparam signed [DEBIT:0]  W_0_x610 = - 23'd388;
localparam signed [DEBIT:0]  W_0_x611 = - 23'd99;
localparam signed [DEBIT:0]  W_0_x612 =  23'd397;
localparam signed [DEBIT:0]  W_0_x613 =  23'd735;
localparam signed [DEBIT:0]  W_0_x614 =  23'd935;
localparam signed [DEBIT:0]  W_0_x615 =  23'd959;
localparam signed [DEBIT:0]  W_0_x616 =  23'd972;
localparam signed [DEBIT:0]  W_0_x617 =  23'd965;
localparam signed [DEBIT:0]  W_0_x618 =  23'd960;
localparam signed [DEBIT:0]  W_0_x619 =  23'd919;
localparam signed [DEBIT:0]  W_0_x620 =  23'd788;
localparam signed [DEBIT:0]  W_0_x621 =  23'd497;
localparam signed [DEBIT:0]  W_0_x622 =  23'd294;
localparam signed [DEBIT:0]  W_0_x623 =  23'd76;
localparam signed [DEBIT:0]  W_0_x624 = - 23'd102;
localparam signed [DEBIT:0]  W_0_x625 =  23'd11;
localparam signed [DEBIT:0]  W_0_x626 =  23'd167;
localparam signed [DEBIT:0]  W_0_x627 =  23'd259;
localparam signed [DEBIT:0]  W_0_x628 =  23'd350;
localparam signed [DEBIT:0]  W_0_x629 =  23'd375;
localparam signed [DEBIT:0]  W_0_x630 =  23'd283;
localparam signed [DEBIT:0]  W_0_x631 =  23'd97;
localparam signed [DEBIT:0]  W_0_x632 =  23'd20;
localparam signed [DEBIT:0]  W_0_x633 = - 23'd80;
localparam signed [DEBIT:0]  W_0_x634 = - 23'd88;
localparam signed [DEBIT:0]  W_0_x635 = - 23'd238;
localparam signed [DEBIT:0]  W_0_x636 = - 23'd326;
localparam signed [DEBIT:0]  W_0_x637 = - 23'd277;
localparam signed [DEBIT:0]  W_0_x638 = - 23'd81;
localparam signed [DEBIT:0]  W_0_x639 =  23'd270;
localparam signed [DEBIT:0]  W_0_x640 =  23'd677;
localparam signed [DEBIT:0]  W_0_x641 =  23'd877;
localparam signed [DEBIT:0]  W_0_x642 =  23'd957;
localparam signed [DEBIT:0]  W_0_x643 =  23'd989;
localparam signed [DEBIT:0]  W_0_x644 =  23'd970;
localparam signed [DEBIT:0]  W_0_x645 =  23'd964;
localparam signed [DEBIT:0]  W_0_x646 =  23'd963;
localparam signed [DEBIT:0]  W_0_x647 =  23'd943;
localparam signed [DEBIT:0]  W_0_x648 =  23'd900;
localparam signed [DEBIT:0]  W_0_x649 =  23'd749;
localparam signed [DEBIT:0]  W_0_x650 =  23'd588;
localparam signed [DEBIT:0]  W_0_x651 =  23'd332;
localparam signed [DEBIT:0]  W_0_x652 =  23'd137;
localparam signed [DEBIT:0]  W_0_x653 =  23'd105;
localparam signed [DEBIT:0]  W_0_x654 =  23'd170;
localparam signed [DEBIT:0]  W_0_x655 =  23'd258;
localparam signed [DEBIT:0]  W_0_x656 =  23'd394;
localparam signed [DEBIT:0]  W_0_x657 =  23'd415;
localparam signed [DEBIT:0]  W_0_x658 =  23'd277;
localparam signed [DEBIT:0]  W_0_x659 =  23'd123;
localparam signed [DEBIT:0]  W_0_x660 =  23'd102;
localparam signed [DEBIT:0]  W_0_x661 =  23'd10;
localparam signed [DEBIT:0]  W_0_x662 = - 23'd23;
localparam signed [DEBIT:0]  W_0_x663 = - 23'd117;
localparam signed [DEBIT:0]  W_0_x664 = - 23'd21;
localparam signed [DEBIT:0]  W_0_x665 =  23'd46;
localparam signed [DEBIT:0]  W_0_x666 =  23'd312;
localparam signed [DEBIT:0]  W_0_x667 =  23'd625;
localparam signed [DEBIT:0]  W_0_x668 =  23'd825;
localparam signed [DEBIT:0]  W_0_x669 =  23'd929;
localparam signed [DEBIT:0]  W_0_x670 =  23'd961;
localparam signed [DEBIT:0]  W_0_x671 =  23'd961;
localparam signed [DEBIT:0]  W_0_x672 =  23'd975;
localparam signed [DEBIT:0]  W_0_x673 =  23'd961;
localparam signed [DEBIT:0]  W_0_x674 =  23'd968;
localparam signed [DEBIT:0]  W_0_x675 =  23'd960;
localparam signed [DEBIT:0]  W_0_x676 =  23'd941;
localparam signed [DEBIT:0]  W_0_x677 =  23'd883;
localparam signed [DEBIT:0]  W_0_x678 =  23'd774;
localparam signed [DEBIT:0]  W_0_x679 =  23'd650;
localparam signed [DEBIT:0]  W_0_x680 =  23'd437;
localparam signed [DEBIT:0]  W_0_x681 =  23'd222;
localparam signed [DEBIT:0]  W_0_x682 = - 23'd28;
localparam signed [DEBIT:0]  W_0_x683 = - 23'd112;
localparam signed [DEBIT:0]  W_0_x684 = - 23'd30;
localparam signed [DEBIT:0]  W_0_x685 =  23'd122;
localparam signed [DEBIT:0]  W_0_x686 =  23'd51;
localparam signed [DEBIT:0]  W_0_x687 =  23'd32;
localparam signed [DEBIT:0]  W_0_x688 =  23'd18;
localparam signed [DEBIT:0]  W_0_x689 =  23'd27;
localparam signed [DEBIT:0]  W_0_x690 =  23'd112;
localparam signed [DEBIT:0]  W_0_x691 =  23'd228;
localparam signed [DEBIT:0]  W_0_x692 =  23'd405;
localparam signed [DEBIT:0]  W_0_x693 =  23'd479;
localparam signed [DEBIT:0]  W_0_x694 =  23'd627;
localparam signed [DEBIT:0]  W_0_x695 =  23'd769;
localparam signed [DEBIT:0]  W_0_x696 =  23'd899;
localparam signed [DEBIT:0]  W_0_x697 =  23'd962;
localparam signed [DEBIT:0]  W_0_x698 =  23'd961;
localparam signed [DEBIT:0]  W_0_x699 =  23'd967;
localparam signed [DEBIT:0]  W_0_x700 =  23'd964;
localparam signed [DEBIT:0]  W_0_x701 =  23'd962;
localparam signed [DEBIT:0]  W_0_x702 =  23'd968;
localparam signed [DEBIT:0]  W_0_x703 =  23'd964;
localparam signed [DEBIT:0]  W_0_x704 =  23'd957;
localparam signed [DEBIT:0]  W_0_x705 =  23'd938;
localparam signed [DEBIT:0]  W_0_x706 =  23'd900;
localparam signed [DEBIT:0]  W_0_x707 =  23'd806;
localparam signed [DEBIT:0]  W_0_x708 =  23'd728;
localparam signed [DEBIT:0]  W_0_x709 =  23'd579;
localparam signed [DEBIT:0]  W_0_x710 =  23'd401;
localparam signed [DEBIT:0]  W_0_x711 =  23'd324;
localparam signed [DEBIT:0]  W_0_x712 =  23'd360;
localparam signed [DEBIT:0]  W_0_x713 =  23'd295;
localparam signed [DEBIT:0]  W_0_x714 =  23'd261;
localparam signed [DEBIT:0]  W_0_x715 =  23'd255;
localparam signed [DEBIT:0]  W_0_x716 =  23'd287;
localparam signed [DEBIT:0]  W_0_x717 =  23'd341;
localparam signed [DEBIT:0]  W_0_x718 =  23'd457;
localparam signed [DEBIT:0]  W_0_x719 =  23'd534;
localparam signed [DEBIT:0]  W_0_x720 =  23'd675;
localparam signed [DEBIT:0]  W_0_x721 =  23'd720;
localparam signed [DEBIT:0]  W_0_x722 =  23'd807;
localparam signed [DEBIT:0]  W_0_x723 =  23'd867;
localparam signed [DEBIT:0]  W_0_x724 =  23'd948;
localparam signed [DEBIT:0]  W_0_x725 =  23'd969;
localparam signed [DEBIT:0]  W_0_x726 =  23'd957;
localparam signed [DEBIT:0]  W_0_x727 =  23'd960;
localparam signed [DEBIT:0]  W_0_x728 =  23'd968;
localparam signed [DEBIT:0]  W_0_x729 =  23'd966;
localparam signed [DEBIT:0]  W_0_x730 =  23'd963;
localparam signed [DEBIT:0]  W_0_x731 =  23'd964;
localparam signed [DEBIT:0]  W_0_x732 =  23'd972;
localparam signed [DEBIT:0]  W_0_x733 =  23'd965;
localparam signed [DEBIT:0]  W_0_x734 =  23'd940;
localparam signed [DEBIT:0]  W_0_x735 =  23'd885;
localparam signed [DEBIT:0]  W_0_x736 =  23'd843;
localparam signed [DEBIT:0]  W_0_x737 =  23'd786;
localparam signed [DEBIT:0]  W_0_x738 =  23'd736;
localparam signed [DEBIT:0]  W_0_x739 =  23'd702;
localparam signed [DEBIT:0]  W_0_x740 =  23'd666;
localparam signed [DEBIT:0]  W_0_x741 =  23'd654;
localparam signed [DEBIT:0]  W_0_x742 =  23'd594;
localparam signed [DEBIT:0]  W_0_x743 =  23'd562;
localparam signed [DEBIT:0]  W_0_x744 =  23'd573;
localparam signed [DEBIT:0]  W_0_x745 =  23'd609;
localparam signed [DEBIT:0]  W_0_x746 =  23'd680;
localparam signed [DEBIT:0]  W_0_x747 =  23'd712;
localparam signed [DEBIT:0]  W_0_x748 =  23'd794;
localparam signed [DEBIT:0]  W_0_x749 =  23'd846;
localparam signed [DEBIT:0]  W_0_x750 =  23'd883;
localparam signed [DEBIT:0]  W_0_x751 =  23'd924;
localparam signed [DEBIT:0]  W_0_x752 =  23'd949;
localparam signed [DEBIT:0]  W_0_x753 =  23'd961;
localparam signed [DEBIT:0]  W_0_x754 =  23'd977;
localparam signed [DEBIT:0]  W_0_x755 =  23'd976;
localparam signed [DEBIT:0]  W_0_x756 =  23'd976;
localparam signed [DEBIT:0]  W_0_x757 =  23'd963;
localparam signed [DEBIT:0]  W_0_x758 =  23'd966;
localparam signed [DEBIT:0]  W_0_x759 =  23'd970;
localparam signed [DEBIT:0]  W_0_x760 =  23'd961;
localparam signed [DEBIT:0]  W_0_x761 =  23'd961;
localparam signed [DEBIT:0]  W_0_x762 =  23'd954;
localparam signed [DEBIT:0]  W_0_x763 =  23'd942;
localparam signed [DEBIT:0]  W_0_x764 =  23'd935;
localparam signed [DEBIT:0]  W_0_x765 =  23'd939;
localparam signed [DEBIT:0]  W_0_x766 =  23'd956;
localparam signed [DEBIT:0]  W_0_x767 =  23'd950;
localparam signed [DEBIT:0]  W_0_x768 =  23'd922;
localparam signed [DEBIT:0]  W_0_x769 =  23'd873;
localparam signed [DEBIT:0]  W_0_x770 =  23'd848;
localparam signed [DEBIT:0]  W_0_x771 =  23'd825;
localparam signed [DEBIT:0]  W_0_x772 =  23'd833;
localparam signed [DEBIT:0]  W_0_x773 =  23'd854;
localparam signed [DEBIT:0]  W_0_x774 =  23'd854;
localparam signed [DEBIT:0]  W_0_x775 =  23'd875;
localparam signed [DEBIT:0]  W_0_x776 =  23'd916;
localparam signed [DEBIT:0]  W_0_x777 =  23'd919;
localparam signed [DEBIT:0]  W_0_x778 =  23'd942;
localparam signed [DEBIT:0]  W_0_x779 =  23'd948;
localparam signed [DEBIT:0]  W_0_x780 =  23'd962;
localparam signed [DEBIT:0]  W_0_x781 =  23'd971;
localparam signed [DEBIT:0]  W_0_x782 =  23'd969;
localparam signed [DEBIT:0]  W_0_x783 =  23'd971;
localparam signed [DEBIT:0]  W_0_x784 =  23'd970;
localparam signed [DEBIT:0]  W_1_x1 =  23'd980;
localparam signed [DEBIT:0]  W_1_x2 =  23'd977;
localparam signed [DEBIT:0]  W_1_x3 =  23'd975;
localparam signed [DEBIT:0]  W_1_x4 =  23'd972;
localparam signed [DEBIT:0]  W_1_x5 =  23'd976;
localparam signed [DEBIT:0]  W_1_x6 =  23'd974;
localparam signed [DEBIT:0]  W_1_x7 =  23'd976;
localparam signed [DEBIT:0]  W_1_x8 =  23'd984;
localparam signed [DEBIT:0]  W_1_x9 =  23'd979;
localparam signed [DEBIT:0]  W_1_x10 =  23'd979;
localparam signed [DEBIT:0]  W_1_x11 =  23'd971;
localparam signed [DEBIT:0]  W_1_x12 =  23'd985;
localparam signed [DEBIT:0]  W_1_x13 =  23'd979;
localparam signed [DEBIT:0]  W_1_x14 =  23'd982;
localparam signed [DEBIT:0]  W_1_x15 =  23'd984;
localparam signed [DEBIT:0]  W_1_x16 =  23'd983;
localparam signed [DEBIT:0]  W_1_x17 =  23'd980;
localparam signed [DEBIT:0]  W_1_x18 =  23'd980;
localparam signed [DEBIT:0]  W_1_x19 =  23'd977;
localparam signed [DEBIT:0]  W_1_x20 =  23'd975;
localparam signed [DEBIT:0]  W_1_x21 =  23'd983;
localparam signed [DEBIT:0]  W_1_x22 =  23'd973;
localparam signed [DEBIT:0]  W_1_x23 =  23'd980;
localparam signed [DEBIT:0]  W_1_x24 =  23'd986;
localparam signed [DEBIT:0]  W_1_x25 =  23'd981;
localparam signed [DEBIT:0]  W_1_x26 =  23'd981;
localparam signed [DEBIT:0]  W_1_x27 =  23'd971;
localparam signed [DEBIT:0]  W_1_x28 =  23'd984;
localparam signed [DEBIT:0]  W_1_x29 =  23'd972;
localparam signed [DEBIT:0]  W_1_x30 =  23'd980;
localparam signed [DEBIT:0]  W_1_x31 =  23'd986;
localparam signed [DEBIT:0]  W_1_x32 =  23'd977;
localparam signed [DEBIT:0]  W_1_x33 =  23'd971;
localparam signed [DEBIT:0]  W_1_x34 =  23'd975;
localparam signed [DEBIT:0]  W_1_x35 =  23'd979;
localparam signed [DEBIT:0]  W_1_x36 =  23'd984;
localparam signed [DEBIT:0]  W_1_x37 =  23'd980;
localparam signed [DEBIT:0]  W_1_x38 =  23'd972;
localparam signed [DEBIT:0]  W_1_x39 =  23'd961;
localparam signed [DEBIT:0]  W_1_x40 =  23'd976;
localparam signed [DEBIT:0]  W_1_x41 =  23'd969;
localparam signed [DEBIT:0]  W_1_x42 =  23'd964;
localparam signed [DEBIT:0]  W_1_x43 =  23'd952;
localparam signed [DEBIT:0]  W_1_x44 =  23'd968;
localparam signed [DEBIT:0]  W_1_x45 =  23'd961;
localparam signed [DEBIT:0]  W_1_x46 =  23'd984;
localparam signed [DEBIT:0]  W_1_x47 =  23'd982;
localparam signed [DEBIT:0]  W_1_x48 =  23'd980;
localparam signed [DEBIT:0]  W_1_x49 =  23'd987;
localparam signed [DEBIT:0]  W_1_x50 =  23'd980;
localparam signed [DEBIT:0]  W_1_x51 =  23'd980;
localparam signed [DEBIT:0]  W_1_x52 =  23'd980;
localparam signed [DEBIT:0]  W_1_x53 =  23'd990;
localparam signed [DEBIT:0]  W_1_x54 =  23'd980;
localparam signed [DEBIT:0]  W_1_x55 =  23'd978;
localparam signed [DEBIT:0]  W_1_x56 =  23'd985;
localparam signed [DEBIT:0]  W_1_x57 =  23'd984;
localparam signed [DEBIT:0]  W_1_x58 =  23'd977;
localparam signed [DEBIT:0]  W_1_x59 =  23'd978;
localparam signed [DEBIT:0]  W_1_x60 =  23'd983;
localparam signed [DEBIT:0]  W_1_x61 =  23'd976;
localparam signed [DEBIT:0]  W_1_x62 =  23'd986;
localparam signed [DEBIT:0]  W_1_x63 =  23'd983;
localparam signed [DEBIT:0]  W_1_x64 =  23'd977;
localparam signed [DEBIT:0]  W_1_x65 =  23'd928;
localparam signed [DEBIT:0]  W_1_x66 =  23'd890;
localparam signed [DEBIT:0]  W_1_x67 =  23'd890;
localparam signed [DEBIT:0]  W_1_x68 =  23'd869;
localparam signed [DEBIT:0]  W_1_x69 =  23'd873;
localparam signed [DEBIT:0]  W_1_x70 =  23'd852;
localparam signed [DEBIT:0]  W_1_x71 =  23'd837;
localparam signed [DEBIT:0]  W_1_x72 =  23'd884;
localparam signed [DEBIT:0]  W_1_x73 =  23'd872;
localparam signed [DEBIT:0]  W_1_x74 =  23'd871;
localparam signed [DEBIT:0]  W_1_x75 =  23'd914;
localparam signed [DEBIT:0]  W_1_x76 =  23'd943;
localparam signed [DEBIT:0]  W_1_x77 =  23'd962;
localparam signed [DEBIT:0]  W_1_x78 =  23'd964;
localparam signed [DEBIT:0]  W_1_x79 =  23'd975;
localparam signed [DEBIT:0]  W_1_x80 =  23'd982;
localparam signed [DEBIT:0]  W_1_x81 =  23'd978;
localparam signed [DEBIT:0]  W_1_x82 =  23'd981;
localparam signed [DEBIT:0]  W_1_x83 =  23'd985;
localparam signed [DEBIT:0]  W_1_x84 =  23'd982;
localparam signed [DEBIT:0]  W_1_x85 =  23'd976;
localparam signed [DEBIT:0]  W_1_x86 =  23'd976;
localparam signed [DEBIT:0]  W_1_x87 =  23'd983;
localparam signed [DEBIT:0]  W_1_x88 =  23'd986;
localparam signed [DEBIT:0]  W_1_x89 =  23'd983;
localparam signed [DEBIT:0]  W_1_x90 =  23'd978;
localparam signed [DEBIT:0]  W_1_x91 =  23'd945;
localparam signed [DEBIT:0]  W_1_x92 =  23'd854;
localparam signed [DEBIT:0]  W_1_x93 =  23'd738;
localparam signed [DEBIT:0]  W_1_x94 =  23'd614;
localparam signed [DEBIT:0]  W_1_x95 =  23'd510;
localparam signed [DEBIT:0]  W_1_x96 =  23'd409;
localparam signed [DEBIT:0]  W_1_x97 =  23'd433;
localparam signed [DEBIT:0]  W_1_x98 =  23'd472;
localparam signed [DEBIT:0]  W_1_x99 =  23'd484;
localparam signed [DEBIT:0]  W_1_x100 =  23'd487;
localparam signed [DEBIT:0]  W_1_x101 =  23'd524;
localparam signed [DEBIT:0]  W_1_x102 =  23'd541;
localparam signed [DEBIT:0]  W_1_x103 =  23'd586;
localparam signed [DEBIT:0]  W_1_x104 =  23'd641;
localparam signed [DEBIT:0]  W_1_x105 =  23'd736;
localparam signed [DEBIT:0]  W_1_x106 =  23'd841;
localparam signed [DEBIT:0]  W_1_x107 =  23'd936;
localparam signed [DEBIT:0]  W_1_x108 =  23'd956;
localparam signed [DEBIT:0]  W_1_x109 =  23'd961;
localparam signed [DEBIT:0]  W_1_x110 =  23'd977;
localparam signed [DEBIT:0]  W_1_x111 =  23'd981;
localparam signed [DEBIT:0]  W_1_x112 =  23'd987;
localparam signed [DEBIT:0]  W_1_x113 =  23'd974;
localparam signed [DEBIT:0]  W_1_x114 =  23'd979;
localparam signed [DEBIT:0]  W_1_x115 =  23'd985;
localparam signed [DEBIT:0]  W_1_x116 =  23'd975;
localparam signed [DEBIT:0]  W_1_x117 =  23'd965;
localparam signed [DEBIT:0]  W_1_x118 =  23'd920;
localparam signed [DEBIT:0]  W_1_x119 =  23'd796;
localparam signed [DEBIT:0]  W_1_x120 =  23'd628;
localparam signed [DEBIT:0]  W_1_x121 =  23'd416;
localparam signed [DEBIT:0]  W_1_x122 =  23'd208;
localparam signed [DEBIT:0]  W_1_x123 =  23'd140;
localparam signed [DEBIT:0]  W_1_x124 =  23'd116;
localparam signed [DEBIT:0]  W_1_x125 =  23'd216;
localparam signed [DEBIT:0]  W_1_x126 =  23'd335;
localparam signed [DEBIT:0]  W_1_x127 =  23'd346;
localparam signed [DEBIT:0]  W_1_x128 =  23'd284;
localparam signed [DEBIT:0]  W_1_x129 =  23'd199;
localparam signed [DEBIT:0]  W_1_x130 =  23'd302;
localparam signed [DEBIT:0]  W_1_x131 =  23'd361;
localparam signed [DEBIT:0]  W_1_x132 =  23'd440;
localparam signed [DEBIT:0]  W_1_x133 =  23'd531;
localparam signed [DEBIT:0]  W_1_x134 =  23'd691;
localparam signed [DEBIT:0]  W_1_x135 =  23'd778;
localparam signed [DEBIT:0]  W_1_x136 =  23'd831;
localparam signed [DEBIT:0]  W_1_x137 =  23'd894;
localparam signed [DEBIT:0]  W_1_x138 =  23'd962;
localparam signed [DEBIT:0]  W_1_x139 =  23'd991;
localparam signed [DEBIT:0]  W_1_x140 =  23'd986;
localparam signed [DEBIT:0]  W_1_x141 =  23'd979;
localparam signed [DEBIT:0]  W_1_x142 =  23'd974;
localparam signed [DEBIT:0]  W_1_x143 =  23'd987;
localparam signed [DEBIT:0]  W_1_x144 =  23'd960;
localparam signed [DEBIT:0]  W_1_x145 =  23'd942;
localparam signed [DEBIT:0]  W_1_x146 =  23'd782;
localparam signed [DEBIT:0]  W_1_x147 =  23'd499;
localparam signed [DEBIT:0]  W_1_x148 =  23'd203;
localparam signed [DEBIT:0]  W_1_x149 = - 23'd84;
localparam signed [DEBIT:0]  W_1_x150 = - 23'd244;
localparam signed [DEBIT:0]  W_1_x151 = - 23'd200;
localparam signed [DEBIT:0]  W_1_x152 = - 23'd153;
localparam signed [DEBIT:0]  W_1_x153 = - 23'd78;
localparam signed [DEBIT:0]  W_1_x154 = - 23'd39;
localparam signed [DEBIT:0]  W_1_x155 =  23'd109;
localparam signed [DEBIT:0]  W_1_x156 =  23'd119;
localparam signed [DEBIT:0]  W_1_x157 =  23'd0;
localparam signed [DEBIT:0]  W_1_x158 =  23'd4;
localparam signed [DEBIT:0]  W_1_x159 =  23'd113;
localparam signed [DEBIT:0]  W_1_x160 =  23'd267;
localparam signed [DEBIT:0]  W_1_x161 =  23'd331;
localparam signed [DEBIT:0]  W_1_x162 =  23'd378;
localparam signed [DEBIT:0]  W_1_x163 =  23'd489;
localparam signed [DEBIT:0]  W_1_x164 =  23'd616;
localparam signed [DEBIT:0]  W_1_x165 =  23'd733;
localparam signed [DEBIT:0]  W_1_x166 =  23'd876;
localparam signed [DEBIT:0]  W_1_x167 =  23'd963;
localparam signed [DEBIT:0]  W_1_x168 =  23'd987;
localparam signed [DEBIT:0]  W_1_x169 =  23'd979;
localparam signed [DEBIT:0]  W_1_x170 =  23'd982;
localparam signed [DEBIT:0]  W_1_x171 =  23'd965;
localparam signed [DEBIT:0]  W_1_x172 =  23'd916;
localparam signed [DEBIT:0]  W_1_x173 =  23'd796;
localparam signed [DEBIT:0]  W_1_x174 =  23'd552;
localparam signed [DEBIT:0]  W_1_x175 =  23'd235;
localparam signed [DEBIT:0]  W_1_x176 = - 23'd80;
localparam signed [DEBIT:0]  W_1_x177 = - 23'd324;
localparam signed [DEBIT:0]  W_1_x178 = - 23'd391;
localparam signed [DEBIT:0]  W_1_x179 = - 23'd337;
localparam signed [DEBIT:0]  W_1_x180 = - 23'd169;
localparam signed [DEBIT:0]  W_1_x181 = - 23'd85;
localparam signed [DEBIT:0]  W_1_x182 = - 23'd91;
localparam signed [DEBIT:0]  W_1_x183 = - 23'd37;
localparam signed [DEBIT:0]  W_1_x184 = - 23'd149;
localparam signed [DEBIT:0]  W_1_x185 = - 23'd112;
localparam signed [DEBIT:0]  W_1_x186 = - 23'd91;
localparam signed [DEBIT:0]  W_1_x187 =  23'd12;
localparam signed [DEBIT:0]  W_1_x188 =  23'd50;
localparam signed [DEBIT:0]  W_1_x189 =  23'd21;
localparam signed [DEBIT:0]  W_1_x190 = - 23'd73;
localparam signed [DEBIT:0]  W_1_x191 =  23'd105;
localparam signed [DEBIT:0]  W_1_x192 =  23'd407;
localparam signed [DEBIT:0]  W_1_x193 =  23'd584;
localparam signed [DEBIT:0]  W_1_x194 =  23'd764;
localparam signed [DEBIT:0]  W_1_x195 =  23'd921;
localparam signed [DEBIT:0]  W_1_x196 =  23'd967;
localparam signed [DEBIT:0]  W_1_x197 =  23'd985;
localparam signed [DEBIT:0]  W_1_x198 =  23'd981;
localparam signed [DEBIT:0]  W_1_x199 =  23'd947;
localparam signed [DEBIT:0]  W_1_x200 =  23'd824;
localparam signed [DEBIT:0]  W_1_x201 =  23'd663;
localparam signed [DEBIT:0]  W_1_x202 =  23'd366;
localparam signed [DEBIT:0]  W_1_x203 =  23'd40;
localparam signed [DEBIT:0]  W_1_x204 = - 23'd189;
localparam signed [DEBIT:0]  W_1_x205 = - 23'd338;
localparam signed [DEBIT:0]  W_1_x206 = - 23'd368;
localparam signed [DEBIT:0]  W_1_x207 = - 23'd225;
localparam signed [DEBIT:0]  W_1_x208 = - 23'd85;
localparam signed [DEBIT:0]  W_1_x209 = - 23'd38;
localparam signed [DEBIT:0]  W_1_x210 = - 23'd116;
localparam signed [DEBIT:0]  W_1_x211 = - 23'd206;
localparam signed [DEBIT:0]  W_1_x212 = - 23'd395;
localparam signed [DEBIT:0]  W_1_x213 = - 23'd363;
localparam signed [DEBIT:0]  W_1_x214 = - 23'd203;
localparam signed [DEBIT:0]  W_1_x215 = - 23'd37;
localparam signed [DEBIT:0]  W_1_x216 =  23'd28;
localparam signed [DEBIT:0]  W_1_x217 = - 23'd123;
localparam signed [DEBIT:0]  W_1_x218 = - 23'd196;
localparam signed [DEBIT:0]  W_1_x219 = - 23'd67;
localparam signed [DEBIT:0]  W_1_x220 =  23'd237;
localparam signed [DEBIT:0]  W_1_x221 =  23'd538;
localparam signed [DEBIT:0]  W_1_x222 =  23'd756;
localparam signed [DEBIT:0]  W_1_x223 =  23'd910;
localparam signed [DEBIT:0]  W_1_x224 =  23'd973;
localparam signed [DEBIT:0]  W_1_x225 =  23'd971;
localparam signed [DEBIT:0]  W_1_x226 =  23'd966;
localparam signed [DEBIT:0]  W_1_x227 =  23'd904;
localparam signed [DEBIT:0]  W_1_x228 =  23'd735;
localparam signed [DEBIT:0]  W_1_x229 =  23'd490;
localparam signed [DEBIT:0]  W_1_x230 =  23'd229;
localparam signed [DEBIT:0]  W_1_x231 = - 23'd111;
localparam signed [DEBIT:0]  W_1_x232 = - 23'd279;
localparam signed [DEBIT:0]  W_1_x233 = - 23'd385;
localparam signed [DEBIT:0]  W_1_x234 = - 23'd349;
localparam signed [DEBIT:0]  W_1_x235 = - 23'd251;
localparam signed [DEBIT:0]  W_1_x236 = - 23'd156;
localparam signed [DEBIT:0]  W_1_x237 = - 23'd123;
localparam signed [DEBIT:0]  W_1_x238 = - 23'd165;
localparam signed [DEBIT:0]  W_1_x239 = - 23'd188;
localparam signed [DEBIT:0]  W_1_x240 = - 23'd259;
localparam signed [DEBIT:0]  W_1_x241 = - 23'd283;
localparam signed [DEBIT:0]  W_1_x242 = - 23'd189;
localparam signed [DEBIT:0]  W_1_x243 = - 23'd137;
localparam signed [DEBIT:0]  W_1_x244 = - 23'd215;
localparam signed [DEBIT:0]  W_1_x245 = - 23'd336;
localparam signed [DEBIT:0]  W_1_x246 = - 23'd381;
localparam signed [DEBIT:0]  W_1_x247 = - 23'd148;
localparam signed [DEBIT:0]  W_1_x248 =  23'd167;
localparam signed [DEBIT:0]  W_1_x249 =  23'd525;
localparam signed [DEBIT:0]  W_1_x250 =  23'd757;
localparam signed [DEBIT:0]  W_1_x251 =  23'd928;
localparam signed [DEBIT:0]  W_1_x252 =  23'd984;
localparam signed [DEBIT:0]  W_1_x253 =  23'd982;
localparam signed [DEBIT:0]  W_1_x254 =  23'd953;
localparam signed [DEBIT:0]  W_1_x255 =  23'd884;
localparam signed [DEBIT:0]  W_1_x256 =  23'd719;
localparam signed [DEBIT:0]  W_1_x257 =  23'd464;
localparam signed [DEBIT:0]  W_1_x258 =  23'd168;
localparam signed [DEBIT:0]  W_1_x259 = - 23'd164;
localparam signed [DEBIT:0]  W_1_x260 = - 23'd287;
localparam signed [DEBIT:0]  W_1_x261 = - 23'd321;
localparam signed [DEBIT:0]  W_1_x262 = - 23'd308;
localparam signed [DEBIT:0]  W_1_x263 = - 23'd238;
localparam signed [DEBIT:0]  W_1_x264 = - 23'd163;
localparam signed [DEBIT:0]  W_1_x265 = - 23'd121;
localparam signed [DEBIT:0]  W_1_x266 = - 23'd125;
localparam signed [DEBIT:0]  W_1_x267 = - 23'd18;
localparam signed [DEBIT:0]  W_1_x268 =  23'd53;
localparam signed [DEBIT:0]  W_1_x269 = - 23'd73;
localparam signed [DEBIT:0]  W_1_x270 = - 23'd265;
localparam signed [DEBIT:0]  W_1_x271 = - 23'd298;
localparam signed [DEBIT:0]  W_1_x272 = - 23'd422;
localparam signed [DEBIT:0]  W_1_x273 = - 23'd487;
localparam signed [DEBIT:0]  W_1_x274 = - 23'd461;
localparam signed [DEBIT:0]  W_1_x275 = - 23'd199;
localparam signed [DEBIT:0]  W_1_x276 =  23'd192;
localparam signed [DEBIT:0]  W_1_x277 =  23'd594;
localparam signed [DEBIT:0]  W_1_x278 =  23'd806;
localparam signed [DEBIT:0]  W_1_x279 =  23'd943;
localparam signed [DEBIT:0]  W_1_x280 =  23'd975;
localparam signed [DEBIT:0]  W_1_x281 =  23'd974;
localparam signed [DEBIT:0]  W_1_x282 =  23'd946;
localparam signed [DEBIT:0]  W_1_x283 =  23'd881;
localparam signed [DEBIT:0]  W_1_x284 =  23'd730;
localparam signed [DEBIT:0]  W_1_x285 =  23'd509;
localparam signed [DEBIT:0]  W_1_x286 =  23'd192;
localparam signed [DEBIT:0]  W_1_x287 = - 23'd156;
localparam signed [DEBIT:0]  W_1_x288 = - 23'd238;
localparam signed [DEBIT:0]  W_1_x289 = - 23'd213;
localparam signed [DEBIT:0]  W_1_x290 = - 23'd136;
localparam signed [DEBIT:0]  W_1_x291 = - 23'd206;
localparam signed [DEBIT:0]  W_1_x292 = - 23'd226;
localparam signed [DEBIT:0]  W_1_x293 = - 23'd103;
localparam signed [DEBIT:0]  W_1_x294 = - 23'd11;
localparam signed [DEBIT:0]  W_1_x295 =  23'd251;
localparam signed [DEBIT:0]  W_1_x296 =  23'd284;
localparam signed [DEBIT:0]  W_1_x297 = - 23'd102;
localparam signed [DEBIT:0]  W_1_x298 = - 23'd298;
localparam signed [DEBIT:0]  W_1_x299 = - 23'd307;
localparam signed [DEBIT:0]  W_1_x300 = - 23'd414;
localparam signed [DEBIT:0]  W_1_x301 = - 23'd537;
localparam signed [DEBIT:0]  W_1_x302 = - 23'd328;
localparam signed [DEBIT:0]  W_1_x303 = - 23'd96;
localparam signed [DEBIT:0]  W_1_x304 =  23'd271;
localparam signed [DEBIT:0]  W_1_x305 =  23'd661;
localparam signed [DEBIT:0]  W_1_x306 =  23'd860;
localparam signed [DEBIT:0]  W_1_x307 =  23'd951;
localparam signed [DEBIT:0]  W_1_x308 =  23'd972;
localparam signed [DEBIT:0]  W_1_x309 =  23'd972;
localparam signed [DEBIT:0]  W_1_x310 =  23'd950;
localparam signed [DEBIT:0]  W_1_x311 =  23'd904;
localparam signed [DEBIT:0]  W_1_x312 =  23'd772;
localparam signed [DEBIT:0]  W_1_x313 =  23'd557;
localparam signed [DEBIT:0]  W_1_x314 =  23'd189;
localparam signed [DEBIT:0]  W_1_x315 = - 23'd197;
localparam signed [DEBIT:0]  W_1_x316 = - 23'd234;
localparam signed [DEBIT:0]  W_1_x317 = - 23'd74;
localparam signed [DEBIT:0]  W_1_x318 = - 23'd51;
localparam signed [DEBIT:0]  W_1_x319 = - 23'd159;
localparam signed [DEBIT:0]  W_1_x320 = - 23'd239;
localparam signed [DEBIT:0]  W_1_x321 = - 23'd186;
localparam signed [DEBIT:0]  W_1_x322 =  23'd49;
localparam signed [DEBIT:0]  W_1_x323 =  23'd399;
localparam signed [DEBIT:0]  W_1_x324 =  23'd391;
localparam signed [DEBIT:0]  W_1_x325 = - 23'd98;
localparam signed [DEBIT:0]  W_1_x326 = - 23'd183;
localparam signed [DEBIT:0]  W_1_x327 = - 23'd184;
localparam signed [DEBIT:0]  W_1_x328 = - 23'd374;
localparam signed [DEBIT:0]  W_1_x329 = - 23'd459;
localparam signed [DEBIT:0]  W_1_x330 = - 23'd213;
localparam signed [DEBIT:0]  W_1_x331 =  23'd17;
localparam signed [DEBIT:0]  W_1_x332 =  23'd350;
localparam signed [DEBIT:0]  W_1_x333 =  23'd676;
localparam signed [DEBIT:0]  W_1_x334 =  23'd896;
localparam signed [DEBIT:0]  W_1_x335 =  23'd962;
localparam signed [DEBIT:0]  W_1_x336 =  23'd976;
localparam signed [DEBIT:0]  W_1_x337 =  23'd984;
localparam signed [DEBIT:0]  W_1_x338 =  23'd956;
localparam signed [DEBIT:0]  W_1_x339 =  23'd912;
localparam signed [DEBIT:0]  W_1_x340 =  23'd834;
localparam signed [DEBIT:0]  W_1_x341 =  23'd603;
localparam signed [DEBIT:0]  W_1_x342 =  23'd172;
localparam signed [DEBIT:0]  W_1_x343 = - 23'd128;
localparam signed [DEBIT:0]  W_1_x344 = - 23'd95;
localparam signed [DEBIT:0]  W_1_x345 =  23'd73;
localparam signed [DEBIT:0]  W_1_x346 = - 23'd5;
localparam signed [DEBIT:0]  W_1_x347 = - 23'd218;
localparam signed [DEBIT:0]  W_1_x348 = - 23'd362;
localparam signed [DEBIT:0]  W_1_x349 = - 23'd276;
localparam signed [DEBIT:0]  W_1_x350 =  23'd174;
localparam signed [DEBIT:0]  W_1_x351 =  23'd607;
localparam signed [DEBIT:0]  W_1_x352 =  23'd397;
localparam signed [DEBIT:0]  W_1_x353 = - 23'd54;
localparam signed [DEBIT:0]  W_1_x354 = - 23'd66;
localparam signed [DEBIT:0]  W_1_x355 = - 23'd127;
localparam signed [DEBIT:0]  W_1_x356 = - 23'd292;
localparam signed [DEBIT:0]  W_1_x357 = - 23'd334;
localparam signed [DEBIT:0]  W_1_x358 = - 23'd111;
localparam signed [DEBIT:0]  W_1_x359 =  23'd78;
localparam signed [DEBIT:0]  W_1_x360 =  23'd363;
localparam signed [DEBIT:0]  W_1_x361 =  23'd651;
localparam signed [DEBIT:0]  W_1_x362 =  23'd895;
localparam signed [DEBIT:0]  W_1_x363 =  23'd969;
localparam signed [DEBIT:0]  W_1_x364 =  23'd979;
localparam signed [DEBIT:0]  W_1_x365 =  23'd982;
localparam signed [DEBIT:0]  W_1_x366 =  23'd969;
localparam signed [DEBIT:0]  W_1_x367 =  23'd948;
localparam signed [DEBIT:0]  W_1_x368 =  23'd877;
localparam signed [DEBIT:0]  W_1_x369 =  23'd676;
localparam signed [DEBIT:0]  W_1_x370 =  23'd254;
localparam signed [DEBIT:0]  W_1_x371 = - 23'd11;
localparam signed [DEBIT:0]  W_1_x372 = - 23'd17;
localparam signed [DEBIT:0]  W_1_x373 =  23'd121;
localparam signed [DEBIT:0]  W_1_x374 = - 23'd13;
localparam signed [DEBIT:0]  W_1_x375 = - 23'd276;
localparam signed [DEBIT:0]  W_1_x376 = - 23'd440;
localparam signed [DEBIT:0]  W_1_x377 = - 23'd254;
localparam signed [DEBIT:0]  W_1_x378 =  23'd267;
localparam signed [DEBIT:0]  W_1_x379 =  23'd562;
localparam signed [DEBIT:0]  W_1_x380 =  23'd270;
localparam signed [DEBIT:0]  W_1_x381 =  23'd47;
localparam signed [DEBIT:0]  W_1_x382 = - 23'd34;
localparam signed [DEBIT:0]  W_1_x383 = - 23'd243;
localparam signed [DEBIT:0]  W_1_x384 = - 23'd234;
localparam signed [DEBIT:0]  W_1_x385 = - 23'd211;
localparam signed [DEBIT:0]  W_1_x386 = - 23'd36;
localparam signed [DEBIT:0]  W_1_x387 =  23'd142;
localparam signed [DEBIT:0]  W_1_x388 =  23'd303;
localparam signed [DEBIT:0]  W_1_x389 =  23'd617;
localparam signed [DEBIT:0]  W_1_x390 =  23'd873;
localparam signed [DEBIT:0]  W_1_x391 =  23'd964;
localparam signed [DEBIT:0]  W_1_x392 =  23'd981;
localparam signed [DEBIT:0]  W_1_x393 =  23'd981;
localparam signed [DEBIT:0]  W_1_x394 =  23'd978;
localparam signed [DEBIT:0]  W_1_x395 =  23'd974;
localparam signed [DEBIT:0]  W_1_x396 =  23'd905;
localparam signed [DEBIT:0]  W_1_x397 =  23'd733;
localparam signed [DEBIT:0]  W_1_x398 =  23'd334;
localparam signed [DEBIT:0]  W_1_x399 =  23'd8;
localparam signed [DEBIT:0]  W_1_x400 = - 23'd43;
localparam signed [DEBIT:0]  W_1_x401 = - 23'd22;
localparam signed [DEBIT:0]  W_1_x402 = - 23'd80;
localparam signed [DEBIT:0]  W_1_x403 = - 23'd331;
localparam signed [DEBIT:0]  W_1_x404 = - 23'd436;
localparam signed [DEBIT:0]  W_1_x405 = - 23'd210;
localparam signed [DEBIT:0]  W_1_x406 =  23'd281;
localparam signed [DEBIT:0]  W_1_x407 =  23'd350;
localparam signed [DEBIT:0]  W_1_x408 =  23'd196;
localparam signed [DEBIT:0]  W_1_x409 =  23'd9;
localparam signed [DEBIT:0]  W_1_x410 = - 23'd251;
localparam signed [DEBIT:0]  W_1_x411 = - 23'd321;
localparam signed [DEBIT:0]  W_1_x412 = - 23'd240;
localparam signed [DEBIT:0]  W_1_x413 = - 23'd146;
localparam signed [DEBIT:0]  W_1_x414 = - 23'd9;
localparam signed [DEBIT:0]  W_1_x415 =  23'd192;
localparam signed [DEBIT:0]  W_1_x416 =  23'd292;
localparam signed [DEBIT:0]  W_1_x417 =  23'd584;
localparam signed [DEBIT:0]  W_1_x418 =  23'd879;
localparam signed [DEBIT:0]  W_1_x419 =  23'd968;
localparam signed [DEBIT:0]  W_1_x420 =  23'd985;
localparam signed [DEBIT:0]  W_1_x421 =  23'd978;
localparam signed [DEBIT:0]  W_1_x422 =  23'd974;
localparam signed [DEBIT:0]  W_1_x423 =  23'd973;
localparam signed [DEBIT:0]  W_1_x424 =  23'd912;
localparam signed [DEBIT:0]  W_1_x425 =  23'd764;
localparam signed [DEBIT:0]  W_1_x426 =  23'd335;
localparam signed [DEBIT:0]  W_1_x427 = - 23'd21;
localparam signed [DEBIT:0]  W_1_x428 = - 23'd131;
localparam signed [DEBIT:0]  W_1_x429 = - 23'd137;
localparam signed [DEBIT:0]  W_1_x430 = - 23'd187;
localparam signed [DEBIT:0]  W_1_x431 = - 23'd332;
localparam signed [DEBIT:0]  W_1_x432 = - 23'd269;
localparam signed [DEBIT:0]  W_1_x433 = - 23'd4;
localparam signed [DEBIT:0]  W_1_x434 =  23'd320;
localparam signed [DEBIT:0]  W_1_x435 =  23'd328;
localparam signed [DEBIT:0]  W_1_x436 =  23'd162;
localparam signed [DEBIT:0]  W_1_x437 = - 23'd57;
localparam signed [DEBIT:0]  W_1_x438 = - 23'd335;
localparam signed [DEBIT:0]  W_1_x439 = - 23'd323;
localparam signed [DEBIT:0]  W_1_x440 = - 23'd253;
localparam signed [DEBIT:0]  W_1_x441 = - 23'd169;
localparam signed [DEBIT:0]  W_1_x442 =  23'd2;
localparam signed [DEBIT:0]  W_1_x443 =  23'd123;
localparam signed [DEBIT:0]  W_1_x444 =  23'd247;
localparam signed [DEBIT:0]  W_1_x445 =  23'd528;
localparam signed [DEBIT:0]  W_1_x446 =  23'd857;
localparam signed [DEBIT:0]  W_1_x447 =  23'd934;
localparam signed [DEBIT:0]  W_1_x448 =  23'd990;
localparam signed [DEBIT:0]  W_1_x449 =  23'd976;
localparam signed [DEBIT:0]  W_1_x450 =  23'd973;
localparam signed [DEBIT:0]  W_1_x451 =  23'd970;
localparam signed [DEBIT:0]  W_1_x452 =  23'd905;
localparam signed [DEBIT:0]  W_1_x453 =  23'd767;
localparam signed [DEBIT:0]  W_1_x454 =  23'd328;
localparam signed [DEBIT:0]  W_1_x455 = - 23'd57;
localparam signed [DEBIT:0]  W_1_x456 = - 23'd251;
localparam signed [DEBIT:0]  W_1_x457 = - 23'd275;
localparam signed [DEBIT:0]  W_1_x458 = - 23'd259;
localparam signed [DEBIT:0]  W_1_x459 = - 23'd199;
localparam signed [DEBIT:0]  W_1_x460 = - 23'd120;
localparam signed [DEBIT:0]  W_1_x461 = - 23'd40;
localparam signed [DEBIT:0]  W_1_x462 =  23'd246;
localparam signed [DEBIT:0]  W_1_x463 =  23'd336;
localparam signed [DEBIT:0]  W_1_x464 =  23'd102;
localparam signed [DEBIT:0]  W_1_x465 = - 23'd153;
localparam signed [DEBIT:0]  W_1_x466 = - 23'd355;
localparam signed [DEBIT:0]  W_1_x467 = - 23'd411;
localparam signed [DEBIT:0]  W_1_x468 = - 23'd340;
localparam signed [DEBIT:0]  W_1_x469 = - 23'd213;
localparam signed [DEBIT:0]  W_1_x470 = - 23'd89;
localparam signed [DEBIT:0]  W_1_x471 =  23'd80;
localparam signed [DEBIT:0]  W_1_x472 =  23'd212;
localparam signed [DEBIT:0]  W_1_x473 =  23'd453;
localparam signed [DEBIT:0]  W_1_x474 =  23'd820;
localparam signed [DEBIT:0]  W_1_x475 =  23'd939;
localparam signed [DEBIT:0]  W_1_x476 =  23'd989;
localparam signed [DEBIT:0]  W_1_x477 =  23'd978;
localparam signed [DEBIT:0]  W_1_x478 =  23'd987;
localparam signed [DEBIT:0]  W_1_x479 =  23'd963;
localparam signed [DEBIT:0]  W_1_x480 =  23'd871;
localparam signed [DEBIT:0]  W_1_x481 =  23'd676;
localparam signed [DEBIT:0]  W_1_x482 =  23'd253;
localparam signed [DEBIT:0]  W_1_x483 = - 23'd137;
localparam signed [DEBIT:0]  W_1_x484 = - 23'd321;
localparam signed [DEBIT:0]  W_1_x485 = - 23'd339;
localparam signed [DEBIT:0]  W_1_x486 = - 23'd236;
localparam signed [DEBIT:0]  W_1_x487 =  23'd10;
localparam signed [DEBIT:0]  W_1_x488 = - 23'd25;
localparam signed [DEBIT:0]  W_1_x489 =  23'd91;
localparam signed [DEBIT:0]  W_1_x490 =  23'd280;
localparam signed [DEBIT:0]  W_1_x491 =  23'd250;
localparam signed [DEBIT:0]  W_1_x492 = - 23'd20;
localparam signed [DEBIT:0]  W_1_x493 = - 23'd226;
localparam signed [DEBIT:0]  W_1_x494 = - 23'd343;
localparam signed [DEBIT:0]  W_1_x495 = - 23'd413;
localparam signed [DEBIT:0]  W_1_x496 = - 23'd330;
localparam signed [DEBIT:0]  W_1_x497 = - 23'd345;
localparam signed [DEBIT:0]  W_1_x498 = - 23'd213;
localparam signed [DEBIT:0]  W_1_x499 =  23'd3;
localparam signed [DEBIT:0]  W_1_x500 =  23'd136;
localparam signed [DEBIT:0]  W_1_x501 =  23'd387;
localparam signed [DEBIT:0]  W_1_x502 =  23'd781;
localparam signed [DEBIT:0]  W_1_x503 =  23'd957;
localparam signed [DEBIT:0]  W_1_x504 =  23'd972;
localparam signed [DEBIT:0]  W_1_x505 =  23'd987;
localparam signed [DEBIT:0]  W_1_x506 =  23'd974;
localparam signed [DEBIT:0]  W_1_x507 =  23'd961;
localparam signed [DEBIT:0]  W_1_x508 =  23'd867;
localparam signed [DEBIT:0]  W_1_x509 =  23'd579;
localparam signed [DEBIT:0]  W_1_x510 =  23'd123;
localparam signed [DEBIT:0]  W_1_x511 = - 23'd216;
localparam signed [DEBIT:0]  W_1_x512 = - 23'd333;
localparam signed [DEBIT:0]  W_1_x513 = - 23'd325;
localparam signed [DEBIT:0]  W_1_x514 = - 23'd197;
localparam signed [DEBIT:0]  W_1_x515 = - 23'd58;
localparam signed [DEBIT:0]  W_1_x516 =  23'd56;
localparam signed [DEBIT:0]  W_1_x517 =  23'd152;
localparam signed [DEBIT:0]  W_1_x518 =  23'd296;
localparam signed [DEBIT:0]  W_1_x519 =  23'd81;
localparam signed [DEBIT:0]  W_1_x520 = - 23'd221;
localparam signed [DEBIT:0]  W_1_x521 = - 23'd273;
localparam signed [DEBIT:0]  W_1_x522 = - 23'd322;
localparam signed [DEBIT:0]  W_1_x523 = - 23'd360;
localparam signed [DEBIT:0]  W_1_x524 = - 23'd330;
localparam signed [DEBIT:0]  W_1_x525 = - 23'd324;
localparam signed [DEBIT:0]  W_1_x526 = - 23'd297;
localparam signed [DEBIT:0]  W_1_x527 = - 23'd198;
localparam signed [DEBIT:0]  W_1_x528 =  23'd94;
localparam signed [DEBIT:0]  W_1_x529 =  23'd439;
localparam signed [DEBIT:0]  W_1_x530 =  23'd828;
localparam signed [DEBIT:0]  W_1_x531 =  23'd964;
localparam signed [DEBIT:0]  W_1_x532 =  23'd982;
localparam signed [DEBIT:0]  W_1_x533 =  23'd975;
localparam signed [DEBIT:0]  W_1_x534 =  23'd982;
localparam signed [DEBIT:0]  W_1_x535 =  23'd935;
localparam signed [DEBIT:0]  W_1_x536 =  23'd779;
localparam signed [DEBIT:0]  W_1_x537 =  23'd479;
localparam signed [DEBIT:0]  W_1_x538 =  23'd88;
localparam signed [DEBIT:0]  W_1_x539 = - 23'd273;
localparam signed [DEBIT:0]  W_1_x540 = - 23'd390;
localparam signed [DEBIT:0]  W_1_x541 = - 23'd377;
localparam signed [DEBIT:0]  W_1_x542 = - 23'd203;
localparam signed [DEBIT:0]  W_1_x543 = - 23'd140;
localparam signed [DEBIT:0]  W_1_x544 = - 23'd95;
localparam signed [DEBIT:0]  W_1_x545 =  23'd5;
localparam signed [DEBIT:0]  W_1_x546 =  23'd142;
localparam signed [DEBIT:0]  W_1_x547 = - 23'd87;
localparam signed [DEBIT:0]  W_1_x548 = - 23'd162;
localparam signed [DEBIT:0]  W_1_x549 = - 23'd187;
localparam signed [DEBIT:0]  W_1_x550 = - 23'd229;
localparam signed [DEBIT:0]  W_1_x551 = - 23'd336;
localparam signed [DEBIT:0]  W_1_x552 = - 23'd381;
localparam signed [DEBIT:0]  W_1_x553 = - 23'd380;
localparam signed [DEBIT:0]  W_1_x554 = - 23'd422;
localparam signed [DEBIT:0]  W_1_x555 = - 23'd273;
localparam signed [DEBIT:0]  W_1_x556 =  23'd109;
localparam signed [DEBIT:0]  W_1_x557 =  23'd545;
localparam signed [DEBIT:0]  W_1_x558 =  23'd859;
localparam signed [DEBIT:0]  W_1_x559 =  23'd971;
localparam signed [DEBIT:0]  W_1_x560 =  23'd972;
localparam signed [DEBIT:0]  W_1_x561 =  23'd985;
localparam signed [DEBIT:0]  W_1_x562 =  23'd968;
localparam signed [DEBIT:0]  W_1_x563 =  23'd925;
localparam signed [DEBIT:0]  W_1_x564 =  23'd744;
localparam signed [DEBIT:0]  W_1_x565 =  23'd424;
localparam signed [DEBIT:0]  W_1_x566 =  23'd43;
localparam signed [DEBIT:0]  W_1_x567 = - 23'd246;
localparam signed [DEBIT:0]  W_1_x568 = - 23'd327;
localparam signed [DEBIT:0]  W_1_x569 = - 23'd252;
localparam signed [DEBIT:0]  W_1_x570 = - 23'd96;
localparam signed [DEBIT:0]  W_1_x571 = - 23'd72;
localparam signed [DEBIT:0]  W_1_x572 = - 23'd94;
localparam signed [DEBIT:0]  W_1_x573 = - 23'd114;
localparam signed [DEBIT:0]  W_1_x574 = - 23'd49;
localparam signed [DEBIT:0]  W_1_x575 = - 23'd164;
localparam signed [DEBIT:0]  W_1_x576 = - 23'd170;
localparam signed [DEBIT:0]  W_1_x577 = - 23'd101;
localparam signed [DEBIT:0]  W_1_x578 = - 23'd112;
localparam signed [DEBIT:0]  W_1_x579 = - 23'd245;
localparam signed [DEBIT:0]  W_1_x580 = - 23'd449;
localparam signed [DEBIT:0]  W_1_x581 = - 23'd521;
localparam signed [DEBIT:0]  W_1_x582 = - 23'd403;
localparam signed [DEBIT:0]  W_1_x583 = - 23'd219;
localparam signed [DEBIT:0]  W_1_x584 =  23'd225;
localparam signed [DEBIT:0]  W_1_x585 =  23'd627;
localparam signed [DEBIT:0]  W_1_x586 =  23'd892;
localparam signed [DEBIT:0]  W_1_x587 =  23'd967;
localparam signed [DEBIT:0]  W_1_x588 =  23'd980;
localparam signed [DEBIT:0]  W_1_x589 =  23'd990;
localparam signed [DEBIT:0]  W_1_x590 =  23'd975;
localparam signed [DEBIT:0]  W_1_x591 =  23'd912;
localparam signed [DEBIT:0]  W_1_x592 =  23'd808;
localparam signed [DEBIT:0]  W_1_x593 =  23'd488;
localparam signed [DEBIT:0]  W_1_x594 =  23'd143;
localparam signed [DEBIT:0]  W_1_x595 = - 23'd140;
localparam signed [DEBIT:0]  W_1_x596 = - 23'd270;
localparam signed [DEBIT:0]  W_1_x597 = - 23'd124;
localparam signed [DEBIT:0]  W_1_x598 = - 23'd55;
localparam signed [DEBIT:0]  W_1_x599 = - 23'd49;
localparam signed [DEBIT:0]  W_1_x600 = - 23'd111;
localparam signed [DEBIT:0]  W_1_x601 = - 23'd196;
localparam signed [DEBIT:0]  W_1_x602 = - 23'd175;
localparam signed [DEBIT:0]  W_1_x603 = - 23'd103;
localparam signed [DEBIT:0]  W_1_x604 =  23'd31;
localparam signed [DEBIT:0]  W_1_x605 = - 23'd11;
localparam signed [DEBIT:0]  W_1_x606 = - 23'd75;
localparam signed [DEBIT:0]  W_1_x607 = - 23'd233;
localparam signed [DEBIT:0]  W_1_x608 = - 23'd421;
localparam signed [DEBIT:0]  W_1_x609 = - 23'd490;
localparam signed [DEBIT:0]  W_1_x610 = - 23'd295;
localparam signed [DEBIT:0]  W_1_x611 = - 23'd34;
localparam signed [DEBIT:0]  W_1_x612 =  23'd472;
localparam signed [DEBIT:0]  W_1_x613 =  23'd758;
localparam signed [DEBIT:0]  W_1_x614 =  23'd934;
localparam signed [DEBIT:0]  W_1_x615 =  23'd967;
localparam signed [DEBIT:0]  W_1_x616 =  23'd985;
localparam signed [DEBIT:0]  W_1_x617 =  23'd983;
localparam signed [DEBIT:0]  W_1_x618 =  23'd980;
localparam signed [DEBIT:0]  W_1_x619 =  23'd932;
localparam signed [DEBIT:0]  W_1_x620 =  23'd877;
localparam signed [DEBIT:0]  W_1_x621 =  23'd632;
localparam signed [DEBIT:0]  W_1_x622 =  23'd397;
localparam signed [DEBIT:0]  W_1_x623 =  23'd135;
localparam signed [DEBIT:0]  W_1_x624 = - 23'd44;
localparam signed [DEBIT:0]  W_1_x625 =  23'd9;
localparam signed [DEBIT:0]  W_1_x626 =  23'd84;
localparam signed [DEBIT:0]  W_1_x627 = - 23'd1;
localparam signed [DEBIT:0]  W_1_x628 = - 23'd186;
localparam signed [DEBIT:0]  W_1_x629 = - 23'd264;
localparam signed [DEBIT:0]  W_1_x630 = - 23'd240;
localparam signed [DEBIT:0]  W_1_x631 =  23'd7;
localparam signed [DEBIT:0]  W_1_x632 =  23'd87;
localparam signed [DEBIT:0]  W_1_x633 =  23'd129;
localparam signed [DEBIT:0]  W_1_x634 =  23'd93;
localparam signed [DEBIT:0]  W_1_x635 = - 23'd62;
localparam signed [DEBIT:0]  W_1_x636 = - 23'd213;
localparam signed [DEBIT:0]  W_1_x637 = - 23'd200;
localparam signed [DEBIT:0]  W_1_x638 = - 23'd10;
localparam signed [DEBIT:0]  W_1_x639 =  23'd312;
localparam signed [DEBIT:0]  W_1_x640 =  23'd672;
localparam signed [DEBIT:0]  W_1_x641 =  23'd855;
localparam signed [DEBIT:0]  W_1_x642 =  23'd961;
localparam signed [DEBIT:0]  W_1_x643 =  23'd987;
localparam signed [DEBIT:0]  W_1_x644 =  23'd980;
localparam signed [DEBIT:0]  W_1_x645 =  23'd978;
localparam signed [DEBIT:0]  W_1_x646 =  23'd989;
localparam signed [DEBIT:0]  W_1_x647 =  23'd967;
localparam signed [DEBIT:0]  W_1_x648 =  23'd930;
localparam signed [DEBIT:0]  W_1_x649 =  23'd820;
localparam signed [DEBIT:0]  W_1_x650 =  23'd673;
localparam signed [DEBIT:0]  W_1_x651 =  23'd456;
localparam signed [DEBIT:0]  W_1_x652 =  23'd266;
localparam signed [DEBIT:0]  W_1_x653 =  23'd193;
localparam signed [DEBIT:0]  W_1_x654 =  23'd165;
localparam signed [DEBIT:0]  W_1_x655 =  23'd12;
localparam signed [DEBIT:0]  W_1_x656 =  23'd7;
localparam signed [DEBIT:0]  W_1_x657 =  23'd14;
localparam signed [DEBIT:0]  W_1_x658 = - 23'd56;
localparam signed [DEBIT:0]  W_1_x659 =  23'd27;
localparam signed [DEBIT:0]  W_1_x660 =  23'd209;
localparam signed [DEBIT:0]  W_1_x661 =  23'd282;
localparam signed [DEBIT:0]  W_1_x662 =  23'd249;
localparam signed [DEBIT:0]  W_1_x663 =  23'd138;
localparam signed [DEBIT:0]  W_1_x664 =  23'd183;
localparam signed [DEBIT:0]  W_1_x665 =  23'd243;
localparam signed [DEBIT:0]  W_1_x666 =  23'd425;
localparam signed [DEBIT:0]  W_1_x667 =  23'd644;
localparam signed [DEBIT:0]  W_1_x668 =  23'd808;
localparam signed [DEBIT:0]  W_1_x669 =  23'd930;
localparam signed [DEBIT:0]  W_1_x670 =  23'd969;
localparam signed [DEBIT:0]  W_1_x671 =  23'd974;
localparam signed [DEBIT:0]  W_1_x672 =  23'd972;
localparam signed [DEBIT:0]  W_1_x673 =  23'd988;
localparam signed [DEBIT:0]  W_1_x674 =  23'd984;
localparam signed [DEBIT:0]  W_1_x675 =  23'd975;
localparam signed [DEBIT:0]  W_1_x676 =  23'd951;
localparam signed [DEBIT:0]  W_1_x677 =  23'd906;
localparam signed [DEBIT:0]  W_1_x678 =  23'd816;
localparam signed [DEBIT:0]  W_1_x679 =  23'd744;
localparam signed [DEBIT:0]  W_1_x680 =  23'd554;
localparam signed [DEBIT:0]  W_1_x681 =  23'd366;
localparam signed [DEBIT:0]  W_1_x682 =  23'd214;
localparam signed [DEBIT:0]  W_1_x683 =  23'd120;
localparam signed [DEBIT:0]  W_1_x684 =  23'd131;
localparam signed [DEBIT:0]  W_1_x685 =  23'd167;
localparam signed [DEBIT:0]  W_1_x686 =  23'd49;
localparam signed [DEBIT:0]  W_1_x687 =  23'd58;
localparam signed [DEBIT:0]  W_1_x688 =  23'd127;
localparam signed [DEBIT:0]  W_1_x689 =  23'd152;
localparam signed [DEBIT:0]  W_1_x690 =  23'd260;
localparam signed [DEBIT:0]  W_1_x691 =  23'd390;
localparam signed [DEBIT:0]  W_1_x692 =  23'd530;
localparam signed [DEBIT:0]  W_1_x693 =  23'd604;
localparam signed [DEBIT:0]  W_1_x694 =  23'd718;
localparam signed [DEBIT:0]  W_1_x695 =  23'd825;
localparam signed [DEBIT:0]  W_1_x696 =  23'd924;
localparam signed [DEBIT:0]  W_1_x697 =  23'd971;
localparam signed [DEBIT:0]  W_1_x698 =  23'd975;
localparam signed [DEBIT:0]  W_1_x699 =  23'd978;
localparam signed [DEBIT:0]  W_1_x700 =  23'd977;
localparam signed [DEBIT:0]  W_1_x701 =  23'd981;
localparam signed [DEBIT:0]  W_1_x702 =  23'd985;
localparam signed [DEBIT:0]  W_1_x703 =  23'd972;
localparam signed [DEBIT:0]  W_1_x704 =  23'd983;
localparam signed [DEBIT:0]  W_1_x705 =  23'd954;
localparam signed [DEBIT:0]  W_1_x706 =  23'd919;
localparam signed [DEBIT:0]  W_1_x707 =  23'd875;
localparam signed [DEBIT:0]  W_1_x708 =  23'd786;
localparam signed [DEBIT:0]  W_1_x709 =  23'd704;
localparam signed [DEBIT:0]  W_1_x710 =  23'd575;
localparam signed [DEBIT:0]  W_1_x711 =  23'd504;
localparam signed [DEBIT:0]  W_1_x712 =  23'd552;
localparam signed [DEBIT:0]  W_1_x713 =  23'd538;
localparam signed [DEBIT:0]  W_1_x714 =  23'd424;
localparam signed [DEBIT:0]  W_1_x715 =  23'd444;
localparam signed [DEBIT:0]  W_1_x716 =  23'd449;
localparam signed [DEBIT:0]  W_1_x717 =  23'd496;
localparam signed [DEBIT:0]  W_1_x718 =  23'd603;
localparam signed [DEBIT:0]  W_1_x719 =  23'd653;
localparam signed [DEBIT:0]  W_1_x720 =  23'd763;
localparam signed [DEBIT:0]  W_1_x721 =  23'd809;
localparam signed [DEBIT:0]  W_1_x722 =  23'd882;
localparam signed [DEBIT:0]  W_1_x723 =  23'd905;
localparam signed [DEBIT:0]  W_1_x724 =  23'd958;
localparam signed [DEBIT:0]  W_1_x725 =  23'd976;
localparam signed [DEBIT:0]  W_1_x726 =  23'd979;
localparam signed [DEBIT:0]  W_1_x727 =  23'd978;
localparam signed [DEBIT:0]  W_1_x728 =  23'd990;
localparam signed [DEBIT:0]  W_1_x729 =  23'd981;
localparam signed [DEBIT:0]  W_1_x730 =  23'd976;
localparam signed [DEBIT:0]  W_1_x731 =  23'd973;
localparam signed [DEBIT:0]  W_1_x732 =  23'd990;
localparam signed [DEBIT:0]  W_1_x733 =  23'd976;
localparam signed [DEBIT:0]  W_1_x734 =  23'd964;
localparam signed [DEBIT:0]  W_1_x735 =  23'd924;
localparam signed [DEBIT:0]  W_1_x736 =  23'd892;
localparam signed [DEBIT:0]  W_1_x737 =  23'd869;
localparam signed [DEBIT:0]  W_1_x738 =  23'd849;
localparam signed [DEBIT:0]  W_1_x739 =  23'd840;
localparam signed [DEBIT:0]  W_1_x740 =  23'd849;
localparam signed [DEBIT:0]  W_1_x741 =  23'd830;
localparam signed [DEBIT:0]  W_1_x742 =  23'd762;
localparam signed [DEBIT:0]  W_1_x743 =  23'd745;
localparam signed [DEBIT:0]  W_1_x744 =  23'd739;
localparam signed [DEBIT:0]  W_1_x745 =  23'd736;
localparam signed [DEBIT:0]  W_1_x746 =  23'd754;
localparam signed [DEBIT:0]  W_1_x747 =  23'd779;
localparam signed [DEBIT:0]  W_1_x748 =  23'd845;
localparam signed [DEBIT:0]  W_1_x749 =  23'd895;
localparam signed [DEBIT:0]  W_1_x750 =  23'd912;
localparam signed [DEBIT:0]  W_1_x751 =  23'd940;
localparam signed [DEBIT:0]  W_1_x752 =  23'd973;
localparam signed [DEBIT:0]  W_1_x753 =  23'd979;
localparam signed [DEBIT:0]  W_1_x754 =  23'd964;
localparam signed [DEBIT:0]  W_1_x755 =  23'd979;
localparam signed [DEBIT:0]  W_1_x756 =  23'd978;
localparam signed [DEBIT:0]  W_1_x757 =  23'd983;
localparam signed [DEBIT:0]  W_1_x758 =  23'd975;
localparam signed [DEBIT:0]  W_1_x759 =  23'd991;
localparam signed [DEBIT:0]  W_1_x760 =  23'd979;
localparam signed [DEBIT:0]  W_1_x761 =  23'd977;
localparam signed [DEBIT:0]  W_1_x762 =  23'd968;
localparam signed [DEBIT:0]  W_1_x763 =  23'd963;
localparam signed [DEBIT:0]  W_1_x764 =  23'd947;
localparam signed [DEBIT:0]  W_1_x765 =  23'd960;
localparam signed [DEBIT:0]  W_1_x766 =  23'd977;
localparam signed [DEBIT:0]  W_1_x767 =  23'd985;
localparam signed [DEBIT:0]  W_1_x768 =  23'd958;
localparam signed [DEBIT:0]  W_1_x769 =  23'd954;
localparam signed [DEBIT:0]  W_1_x770 =  23'd969;
localparam signed [DEBIT:0]  W_1_x771 =  23'd967;
localparam signed [DEBIT:0]  W_1_x772 =  23'd928;
localparam signed [DEBIT:0]  W_1_x773 =  23'd903;
localparam signed [DEBIT:0]  W_1_x774 =  23'd891;
localparam signed [DEBIT:0]  W_1_x775 =  23'd900;
localparam signed [DEBIT:0]  W_1_x776 =  23'd943;
localparam signed [DEBIT:0]  W_1_x777 =  23'd955;
localparam signed [DEBIT:0]  W_1_x778 =  23'd961;
localparam signed [DEBIT:0]  W_1_x779 =  23'd972;
localparam signed [DEBIT:0]  W_1_x780 =  23'd976;
localparam signed [DEBIT:0]  W_1_x781 =  23'd973;
localparam signed [DEBIT:0]  W_1_x782 =  23'd976;
localparam signed [DEBIT:0]  W_1_x783 =  23'd977;
localparam signed [DEBIT:0]  W_1_x784 =  23'd978;
localparam signed [DEBIT:0]  W_2_x1 =  23'd967;
localparam signed [DEBIT:0]  W_2_x2 =  23'd966;
localparam signed [DEBIT:0]  W_2_x3 =  23'd967;
localparam signed [DEBIT:0]  W_2_x4 =  23'd961;
localparam signed [DEBIT:0]  W_2_x5 =  23'd970;
localparam signed [DEBIT:0]  W_2_x6 =  23'd976;
localparam signed [DEBIT:0]  W_2_x7 =  23'd969;
localparam signed [DEBIT:0]  W_2_x8 =  23'd974;
localparam signed [DEBIT:0]  W_2_x9 =  23'd966;
localparam signed [DEBIT:0]  W_2_x10 =  23'd963;
localparam signed [DEBIT:0]  W_2_x11 =  23'd967;
localparam signed [DEBIT:0]  W_2_x12 =  23'd970;
localparam signed [DEBIT:0]  W_2_x13 =  23'd967;
localparam signed [DEBIT:0]  W_2_x14 =  23'd964;
localparam signed [DEBIT:0]  W_2_x15 =  23'd964;
localparam signed [DEBIT:0]  W_2_x16 =  23'd961;
localparam signed [DEBIT:0]  W_2_x17 =  23'd972;
localparam signed [DEBIT:0]  W_2_x18 =  23'd967;
localparam signed [DEBIT:0]  W_2_x19 =  23'd965;
localparam signed [DEBIT:0]  W_2_x20 =  23'd974;
localparam signed [DEBIT:0]  W_2_x21 =  23'd966;
localparam signed [DEBIT:0]  W_2_x22 =  23'd964;
localparam signed [DEBIT:0]  W_2_x23 =  23'd961;
localparam signed [DEBIT:0]  W_2_x24 =  23'd960;
localparam signed [DEBIT:0]  W_2_x25 =  23'd963;
localparam signed [DEBIT:0]  W_2_x26 =  23'd972;
localparam signed [DEBIT:0]  W_2_x27 =  23'd969;
localparam signed [DEBIT:0]  W_2_x28 =  23'd972;
localparam signed [DEBIT:0]  W_2_x29 =  23'd970;
localparam signed [DEBIT:0]  W_2_x30 =  23'd961;
localparam signed [DEBIT:0]  W_2_x31 =  23'd962;
localparam signed [DEBIT:0]  W_2_x32 =  23'd959;
localparam signed [DEBIT:0]  W_2_x33 =  23'd953;
localparam signed [DEBIT:0]  W_2_x34 =  23'd965;
localparam signed [DEBIT:0]  W_2_x35 =  23'd957;
localparam signed [DEBIT:0]  W_2_x36 =  23'd960;
localparam signed [DEBIT:0]  W_2_x37 =  23'd944;
localparam signed [DEBIT:0]  W_2_x38 =  23'd939;
localparam signed [DEBIT:0]  W_2_x39 =  23'd945;
localparam signed [DEBIT:0]  W_2_x40 =  23'd937;
localparam signed [DEBIT:0]  W_2_x41 =  23'd930;
localparam signed [DEBIT:0]  W_2_x42 =  23'd897;
localparam signed [DEBIT:0]  W_2_x43 =  23'd877;
localparam signed [DEBIT:0]  W_2_x44 =  23'd917;
localparam signed [DEBIT:0]  W_2_x45 =  23'd936;
localparam signed [DEBIT:0]  W_2_x46 =  23'd921;
localparam signed [DEBIT:0]  W_2_x47 =  23'd929;
localparam signed [DEBIT:0]  W_2_x48 =  23'd938;
localparam signed [DEBIT:0]  W_2_x49 =  23'd958;
localparam signed [DEBIT:0]  W_2_x50 =  23'd956;
localparam signed [DEBIT:0]  W_2_x51 =  23'd962;
localparam signed [DEBIT:0]  W_2_x52 =  23'd959;
localparam signed [DEBIT:0]  W_2_x53 =  23'd965;
localparam signed [DEBIT:0]  W_2_x54 =  23'd968;
localparam signed [DEBIT:0]  W_2_x55 =  23'd967;
localparam signed [DEBIT:0]  W_2_x56 =  23'd963;
localparam signed [DEBIT:0]  W_2_x57 =  23'd960;
localparam signed [DEBIT:0]  W_2_x58 =  23'd959;
localparam signed [DEBIT:0]  W_2_x59 =  23'd957;
localparam signed [DEBIT:0]  W_2_x60 =  23'd968;
localparam signed [DEBIT:0]  W_2_x61 =  23'd971;
localparam signed [DEBIT:0]  W_2_x62 =  23'd966;
localparam signed [DEBIT:0]  W_2_x63 =  23'd960;
localparam signed [DEBIT:0]  W_2_x64 =  23'd950;
localparam signed [DEBIT:0]  W_2_x65 =  23'd899;
localparam signed [DEBIT:0]  W_2_x66 =  23'd845;
localparam signed [DEBIT:0]  W_2_x67 =  23'd819;
localparam signed [DEBIT:0]  W_2_x68 =  23'd804;
localparam signed [DEBIT:0]  W_2_x69 =  23'd713;
localparam signed [DEBIT:0]  W_2_x70 =  23'd619;
localparam signed [DEBIT:0]  W_2_x71 =  23'd497;
localparam signed [DEBIT:0]  W_2_x72 =  23'd462;
localparam signed [DEBIT:0]  W_2_x73 =  23'd469;
localparam signed [DEBIT:0]  W_2_x74 =  23'd509;
localparam signed [DEBIT:0]  W_2_x75 =  23'd611;
localparam signed [DEBIT:0]  W_2_x76 =  23'd716;
localparam signed [DEBIT:0]  W_2_x77 =  23'd836;
localparam signed [DEBIT:0]  W_2_x78 =  23'd870;
localparam signed [DEBIT:0]  W_2_x79 =  23'd899;
localparam signed [DEBIT:0]  W_2_x80 =  23'd946;
localparam signed [DEBIT:0]  W_2_x81 =  23'd952;
localparam signed [DEBIT:0]  W_2_x82 =  23'd965;
localparam signed [DEBIT:0]  W_2_x83 =  23'd964;
localparam signed [DEBIT:0]  W_2_x84 =  23'd977;
localparam signed [DEBIT:0]  W_2_x85 =  23'd973;
localparam signed [DEBIT:0]  W_2_x86 =  23'd963;
localparam signed [DEBIT:0]  W_2_x87 =  23'd960;
localparam signed [DEBIT:0]  W_2_x88 =  23'd962;
localparam signed [DEBIT:0]  W_2_x89 =  23'd970;
localparam signed [DEBIT:0]  W_2_x90 =  23'd949;
localparam signed [DEBIT:0]  W_2_x91 =  23'd917;
localparam signed [DEBIT:0]  W_2_x92 =  23'd883;
localparam signed [DEBIT:0]  W_2_x93 =  23'd825;
localparam signed [DEBIT:0]  W_2_x94 =  23'd801;
localparam signed [DEBIT:0]  W_2_x95 =  23'd738;
localparam signed [DEBIT:0]  W_2_x96 =  23'd625;
localparam signed [DEBIT:0]  W_2_x97 =  23'd506;
localparam signed [DEBIT:0]  W_2_x98 =  23'd410;
localparam signed [DEBIT:0]  W_2_x99 =  23'd159;
localparam signed [DEBIT:0]  W_2_x100 =  23'd32;
localparam signed [DEBIT:0]  W_2_x101 =  23'd56;
localparam signed [DEBIT:0]  W_2_x102 =  23'd74;
localparam signed [DEBIT:0]  W_2_x103 =  23'd210;
localparam signed [DEBIT:0]  W_2_x104 =  23'd321;
localparam signed [DEBIT:0]  W_2_x105 =  23'd494;
localparam signed [DEBIT:0]  W_2_x106 =  23'd599;
localparam signed [DEBIT:0]  W_2_x107 =  23'd758;
localparam signed [DEBIT:0]  W_2_x108 =  23'd888;
localparam signed [DEBIT:0]  W_2_x109 =  23'd933;
localparam signed [DEBIT:0]  W_2_x110 =  23'd955;
localparam signed [DEBIT:0]  W_2_x111 =  23'd962;
localparam signed [DEBIT:0]  W_2_x112 =  23'd976;
localparam signed [DEBIT:0]  W_2_x113 =  23'd956;
localparam signed [DEBIT:0]  W_2_x114 =  23'd971;
localparam signed [DEBIT:0]  W_2_x115 =  23'd968;
localparam signed [DEBIT:0]  W_2_x116 =  23'd967;
localparam signed [DEBIT:0]  W_2_x117 =  23'd942;
localparam signed [DEBIT:0]  W_2_x118 =  23'd896;
localparam signed [DEBIT:0]  W_2_x119 =  23'd822;
localparam signed [DEBIT:0]  W_2_x120 =  23'd710;
localparam signed [DEBIT:0]  W_2_x121 =  23'd555;
localparam signed [DEBIT:0]  W_2_x122 =  23'd481;
localparam signed [DEBIT:0]  W_2_x123 =  23'd436;
localparam signed [DEBIT:0]  W_2_x124 =  23'd418;
localparam signed [DEBIT:0]  W_2_x125 =  23'd383;
localparam signed [DEBIT:0]  W_2_x126 =  23'd327;
localparam signed [DEBIT:0]  W_2_x127 =  23'd340;
localparam signed [DEBIT:0]  W_2_x128 =  23'd319;
localparam signed [DEBIT:0]  W_2_x129 =  23'd219;
localparam signed [DEBIT:0]  W_2_x130 =  23'd84;
localparam signed [DEBIT:0]  W_2_x131 =  23'd37;
localparam signed [DEBIT:0]  W_2_x132 =  23'd68;
localparam signed [DEBIT:0]  W_2_x133 =  23'd99;
localparam signed [DEBIT:0]  W_2_x134 =  23'd217;
localparam signed [DEBIT:0]  W_2_x135 =  23'd362;
localparam signed [DEBIT:0]  W_2_x136 =  23'd623;
localparam signed [DEBIT:0]  W_2_x137 =  23'd812;
localparam signed [DEBIT:0]  W_2_x138 =  23'd935;
localparam signed [DEBIT:0]  W_2_x139 =  23'd966;
localparam signed [DEBIT:0]  W_2_x140 =  23'd963;
localparam signed [DEBIT:0]  W_2_x141 =  23'd962;
localparam signed [DEBIT:0]  W_2_x142 =  23'd966;
localparam signed [DEBIT:0]  W_2_x143 =  23'd965;
localparam signed [DEBIT:0]  W_2_x144 =  23'd952;
localparam signed [DEBIT:0]  W_2_x145 =  23'd849;
localparam signed [DEBIT:0]  W_2_x146 =  23'd703;
localparam signed [DEBIT:0]  W_2_x147 =  23'd504;
localparam signed [DEBIT:0]  W_2_x148 =  23'd356;
localparam signed [DEBIT:0]  W_2_x149 =  23'd256;
localparam signed [DEBIT:0]  W_2_x150 =  23'd201;
localparam signed [DEBIT:0]  W_2_x151 =  23'd251;
localparam signed [DEBIT:0]  W_2_x152 =  23'd278;
localparam signed [DEBIT:0]  W_2_x153 =  23'd212;
localparam signed [DEBIT:0]  W_2_x154 =  23'd183;
localparam signed [DEBIT:0]  W_2_x155 =  23'd430;
localparam signed [DEBIT:0]  W_2_x156 =  23'd426;
localparam signed [DEBIT:0]  W_2_x157 =  23'd351;
localparam signed [DEBIT:0]  W_2_x158 =  23'd246;
localparam signed [DEBIT:0]  W_2_x159 =  23'd69;
localparam signed [DEBIT:0]  W_2_x160 = - 23'd73;
localparam signed [DEBIT:0]  W_2_x161 = - 23'd119;
localparam signed [DEBIT:0]  W_2_x162 = - 23'd119;
localparam signed [DEBIT:0]  W_2_x163 =  23'd129;
localparam signed [DEBIT:0]  W_2_x164 =  23'd395;
localparam signed [DEBIT:0]  W_2_x165 =  23'd653;
localparam signed [DEBIT:0]  W_2_x166 =  23'd871;
localparam signed [DEBIT:0]  W_2_x167 =  23'd956;
localparam signed [DEBIT:0]  W_2_x168 =  23'd961;
localparam signed [DEBIT:0]  W_2_x169 =  23'd963;
localparam signed [DEBIT:0]  W_2_x170 =  23'd968;
localparam signed [DEBIT:0]  W_2_x171 =  23'd949;
localparam signed [DEBIT:0]  W_2_x172 =  23'd856;
localparam signed [DEBIT:0]  W_2_x173 =  23'd652;
localparam signed [DEBIT:0]  W_2_x174 =  23'd447;
localparam signed [DEBIT:0]  W_2_x175 =  23'd251;
localparam signed [DEBIT:0]  W_2_x176 =  23'd145;
localparam signed [DEBIT:0]  W_2_x177 =  23'd80;
localparam signed [DEBIT:0]  W_2_x178 =  23'd114;
localparam signed [DEBIT:0]  W_2_x179 =  23'd178;
localparam signed [DEBIT:0]  W_2_x180 =  23'd177;
localparam signed [DEBIT:0]  W_2_x181 =  23'd186;
localparam signed [DEBIT:0]  W_2_x182 =  23'd146;
localparam signed [DEBIT:0]  W_2_x183 =  23'd193;
localparam signed [DEBIT:0]  W_2_x184 =  23'd207;
localparam signed [DEBIT:0]  W_2_x185 =  23'd260;
localparam signed [DEBIT:0]  W_2_x186 =  23'd283;
localparam signed [DEBIT:0]  W_2_x187 =  23'd111;
localparam signed [DEBIT:0]  W_2_x188 = - 23'd43;
localparam signed [DEBIT:0]  W_2_x189 = - 23'd245;
localparam signed [DEBIT:0]  W_2_x190 = - 23'd271;
localparam signed [DEBIT:0]  W_2_x191 = - 23'd83;
localparam signed [DEBIT:0]  W_2_x192 =  23'd286;
localparam signed [DEBIT:0]  W_2_x193 =  23'd568;
localparam signed [DEBIT:0]  W_2_x194 =  23'd786;
localparam signed [DEBIT:0]  W_2_x195 =  23'd918;
localparam signed [DEBIT:0]  W_2_x196 =  23'd958;
localparam signed [DEBIT:0]  W_2_x197 =  23'd968;
localparam signed [DEBIT:0]  W_2_x198 =  23'd956;
localparam signed [DEBIT:0]  W_2_x199 =  23'd923;
localparam signed [DEBIT:0]  W_2_x200 =  23'd751;
localparam signed [DEBIT:0]  W_2_x201 =  23'd479;
localparam signed [DEBIT:0]  W_2_x202 =  23'd188;
localparam signed [DEBIT:0]  W_2_x203 =  23'd76;
localparam signed [DEBIT:0]  W_2_x204 = - 23'd69;
localparam signed [DEBIT:0]  W_2_x205 =  23'd16;
localparam signed [DEBIT:0]  W_2_x206 = - 23'd7;
localparam signed [DEBIT:0]  W_2_x207 =  23'd122;
localparam signed [DEBIT:0]  W_2_x208 =  23'd124;
localparam signed [DEBIT:0]  W_2_x209 =  23'd93;
localparam signed [DEBIT:0]  W_2_x210 =  23'd78;
localparam signed [DEBIT:0]  W_2_x211 =  23'd53;
localparam signed [DEBIT:0]  W_2_x212 = - 23'd79;
localparam signed [DEBIT:0]  W_2_x213 = - 23'd59;
localparam signed [DEBIT:0]  W_2_x214 = - 23'd22;
localparam signed [DEBIT:0]  W_2_x215 = - 23'd38;
localparam signed [DEBIT:0]  W_2_x216 = - 23'd7;
localparam signed [DEBIT:0]  W_2_x217 = - 23'd179;
localparam signed [DEBIT:0]  W_2_x218 = - 23'd217;
localparam signed [DEBIT:0]  W_2_x219 = - 23'd66;
localparam signed [DEBIT:0]  W_2_x220 =  23'd184;
localparam signed [DEBIT:0]  W_2_x221 =  23'd496;
localparam signed [DEBIT:0]  W_2_x222 =  23'd741;
localparam signed [DEBIT:0]  W_2_x223 =  23'd888;
localparam signed [DEBIT:0]  W_2_x224 =  23'd957;
localparam signed [DEBIT:0]  W_2_x225 =  23'd965;
localparam signed [DEBIT:0]  W_2_x226 =  23'd925;
localparam signed [DEBIT:0]  W_2_x227 =  23'd836;
localparam signed [DEBIT:0]  W_2_x228 =  23'd578;
localparam signed [DEBIT:0]  W_2_x229 =  23'd270;
localparam signed [DEBIT:0]  W_2_x230 =  23'd82;
localparam signed [DEBIT:0]  W_2_x231 = - 23'd76;
localparam signed [DEBIT:0]  W_2_x232 = - 23'd128;
localparam signed [DEBIT:0]  W_2_x233 = - 23'd127;
localparam signed [DEBIT:0]  W_2_x234 = - 23'd8;
localparam signed [DEBIT:0]  W_2_x235 =  23'd107;
localparam signed [DEBIT:0]  W_2_x236 =  23'd156;
localparam signed [DEBIT:0]  W_2_x237 = - 23'd8;
localparam signed [DEBIT:0]  W_2_x238 = - 23'd24;
localparam signed [DEBIT:0]  W_2_x239 =  23'd0;
localparam signed [DEBIT:0]  W_2_x240 = - 23'd134;
localparam signed [DEBIT:0]  W_2_x241 = - 23'd237;
localparam signed [DEBIT:0]  W_2_x242 = - 23'd151;
localparam signed [DEBIT:0]  W_2_x243 = - 23'd225;
localparam signed [DEBIT:0]  W_2_x244 = - 23'd108;
localparam signed [DEBIT:0]  W_2_x245 = - 23'd155;
localparam signed [DEBIT:0]  W_2_x246 = - 23'd299;
localparam signed [DEBIT:0]  W_2_x247 = - 23'd132;
localparam signed [DEBIT:0]  W_2_x248 =  23'd139;
localparam signed [DEBIT:0]  W_2_x249 =  23'd422;
localparam signed [DEBIT:0]  W_2_x250 =  23'd699;
localparam signed [DEBIT:0]  W_2_x251 =  23'd903;
localparam signed [DEBIT:0]  W_2_x252 =  23'd973;
localparam signed [DEBIT:0]  W_2_x253 =  23'd980;
localparam signed [DEBIT:0]  W_2_x254 =  23'd904;
localparam signed [DEBIT:0]  W_2_x255 =  23'd776;
localparam signed [DEBIT:0]  W_2_x256 =  23'd554;
localparam signed [DEBIT:0]  W_2_x257 =  23'd301;
localparam signed [DEBIT:0]  W_2_x258 =  23'd153;
localparam signed [DEBIT:0]  W_2_x259 = - 23'd74;
localparam signed [DEBIT:0]  W_2_x260 = - 23'd138;
localparam signed [DEBIT:0]  W_2_x261 = - 23'd209;
localparam signed [DEBIT:0]  W_2_x262 = - 23'd70;
localparam signed [DEBIT:0]  W_2_x263 =  23'd47;
localparam signed [DEBIT:0]  W_2_x264 =  23'd108;
localparam signed [DEBIT:0]  W_2_x265 =  23'd9;
localparam signed [DEBIT:0]  W_2_x266 = - 23'd64;
localparam signed [DEBIT:0]  W_2_x267 = - 23'd111;
localparam signed [DEBIT:0]  W_2_x268 = - 23'd26;
localparam signed [DEBIT:0]  W_2_x269 = - 23'd41;
localparam signed [DEBIT:0]  W_2_x270 = - 23'd61;
localparam signed [DEBIT:0]  W_2_x271 = - 23'd132;
localparam signed [DEBIT:0]  W_2_x272 = - 23'd227;
localparam signed [DEBIT:0]  W_2_x273 = - 23'd209;
localparam signed [DEBIT:0]  W_2_x274 = - 23'd329;
localparam signed [DEBIT:0]  W_2_x275 = - 23'd203;
localparam signed [DEBIT:0]  W_2_x276 =  23'd84;
localparam signed [DEBIT:0]  W_2_x277 =  23'd465;
localparam signed [DEBIT:0]  W_2_x278 =  23'd778;
localparam signed [DEBIT:0]  W_2_x279 =  23'd916;
localparam signed [DEBIT:0]  W_2_x280 =  23'd951;
localparam signed [DEBIT:0]  W_2_x281 =  23'd964;
localparam signed [DEBIT:0]  W_2_x282 =  23'd893;
localparam signed [DEBIT:0]  W_2_x283 =  23'd809;
localparam signed [DEBIT:0]  W_2_x284 =  23'd618;
localparam signed [DEBIT:0]  W_2_x285 =  23'd384;
localparam signed [DEBIT:0]  W_2_x286 =  23'd121;
localparam signed [DEBIT:0]  W_2_x287 = - 23'd169;
localparam signed [DEBIT:0]  W_2_x288 = - 23'd267;
localparam signed [DEBIT:0]  W_2_x289 = - 23'd147;
localparam signed [DEBIT:0]  W_2_x290 = - 23'd114;
localparam signed [DEBIT:0]  W_2_x291 = - 23'd141;
localparam signed [DEBIT:0]  W_2_x292 = - 23'd149;
localparam signed [DEBIT:0]  W_2_x293 = - 23'd251;
localparam signed [DEBIT:0]  W_2_x294 = - 23'd304;
localparam signed [DEBIT:0]  W_2_x295 = - 23'd204;
localparam signed [DEBIT:0]  W_2_x296 = - 23'd163;
localparam signed [DEBIT:0]  W_2_x297 = - 23'd199;
localparam signed [DEBIT:0]  W_2_x298 = - 23'd50;
localparam signed [DEBIT:0]  W_2_x299 = - 23'd92;
localparam signed [DEBIT:0]  W_2_x300 = - 23'd115;
localparam signed [DEBIT:0]  W_2_x301 = - 23'd77;
localparam signed [DEBIT:0]  W_2_x302 = - 23'd199;
localparam signed [DEBIT:0]  W_2_x303 = - 23'd209;
localparam signed [DEBIT:0]  W_2_x304 =  23'd69;
localparam signed [DEBIT:0]  W_2_x305 =  23'd549;
localparam signed [DEBIT:0]  W_2_x306 =  23'd833;
localparam signed [DEBIT:0]  W_2_x307 =  23'd933;
localparam signed [DEBIT:0]  W_2_x308 =  23'd957;
localparam signed [DEBIT:0]  W_2_x309 =  23'd966;
localparam signed [DEBIT:0]  W_2_x310 =  23'd913;
localparam signed [DEBIT:0]  W_2_x311 =  23'd858;
localparam signed [DEBIT:0]  W_2_x312 =  23'd705;
localparam signed [DEBIT:0]  W_2_x313 =  23'd455;
localparam signed [DEBIT:0]  W_2_x314 =  23'd49;
localparam signed [DEBIT:0]  W_2_x315 = - 23'd418;
localparam signed [DEBIT:0]  W_2_x316 = - 23'd521;
localparam signed [DEBIT:0]  W_2_x317 = - 23'd336;
localparam signed [DEBIT:0]  W_2_x318 = - 23'd330;
localparam signed [DEBIT:0]  W_2_x319 = - 23'd449;
localparam signed [DEBIT:0]  W_2_x320 = - 23'd491;
localparam signed [DEBIT:0]  W_2_x321 = - 23'd563;
localparam signed [DEBIT:0]  W_2_x322 = - 23'd638;
localparam signed [DEBIT:0]  W_2_x323 = - 23'd591;
localparam signed [DEBIT:0]  W_2_x324 = - 23'd322;
localparam signed [DEBIT:0]  W_2_x325 = - 23'd152;
localparam signed [DEBIT:0]  W_2_x326 = - 23'd6;
localparam signed [DEBIT:0]  W_2_x327 = - 23'd72;
localparam signed [DEBIT:0]  W_2_x328 =  23'd109;
localparam signed [DEBIT:0]  W_2_x329 = - 23'd16;
localparam signed [DEBIT:0]  W_2_x330 = - 23'd213;
localparam signed [DEBIT:0]  W_2_x331 = - 23'd306;
localparam signed [DEBIT:0]  W_2_x332 = - 23'd6;
localparam signed [DEBIT:0]  W_2_x333 =  23'd532;
localparam signed [DEBIT:0]  W_2_x334 =  23'd894;
localparam signed [DEBIT:0]  W_2_x335 =  23'd944;
localparam signed [DEBIT:0]  W_2_x336 =  23'd962;
localparam signed [DEBIT:0]  W_2_x337 =  23'd957;
localparam signed [DEBIT:0]  W_2_x338 =  23'd949;
localparam signed [DEBIT:0]  W_2_x339 =  23'd897;
localparam signed [DEBIT:0]  W_2_x340 =  23'd768;
localparam signed [DEBIT:0]  W_2_x341 =  23'd442;
localparam signed [DEBIT:0]  W_2_x342 = - 23'd152;
localparam signed [DEBIT:0]  W_2_x343 = - 23'd736;
localparam signed [DEBIT:0]  W_2_x344 = - 23'd747;
localparam signed [DEBIT:0]  W_2_x345 = - 23'd523;
localparam signed [DEBIT:0]  W_2_x346 = - 23'd545;
localparam signed [DEBIT:0]  W_2_x347 = - 23'd646;
localparam signed [DEBIT:0]  W_2_x348 = - 23'd726;
localparam signed [DEBIT:0]  W_2_x349 = - 23'd685;
localparam signed [DEBIT:0]  W_2_x350 = - 23'd630;
localparam signed [DEBIT:0]  W_2_x351 = - 23'd624;
localparam signed [DEBIT:0]  W_2_x352 = - 23'd409;
localparam signed [DEBIT:0]  W_2_x353 = - 23'd208;
localparam signed [DEBIT:0]  W_2_x354 = - 23'd250;
localparam signed [DEBIT:0]  W_2_x355 = - 23'd112;
localparam signed [DEBIT:0]  W_2_x356 =  23'd65;
localparam signed [DEBIT:0]  W_2_x357 = - 23'd173;
localparam signed [DEBIT:0]  W_2_x358 = - 23'd246;
localparam signed [DEBIT:0]  W_2_x359 = - 23'd391;
localparam signed [DEBIT:0]  W_2_x360 = - 23'd151;
localparam signed [DEBIT:0]  W_2_x361 =  23'd418;
localparam signed [DEBIT:0]  W_2_x362 =  23'd915;
localparam signed [DEBIT:0]  W_2_x363 =  23'd967;
localparam signed [DEBIT:0]  W_2_x364 =  23'd963;
localparam signed [DEBIT:0]  W_2_x365 =  23'd968;
localparam signed [DEBIT:0]  W_2_x366 =  23'd953;
localparam signed [DEBIT:0]  W_2_x367 =  23'd939;
localparam signed [DEBIT:0]  W_2_x368 =  23'd794;
localparam signed [DEBIT:0]  W_2_x369 =  23'd452;
localparam signed [DEBIT:0]  W_2_x370 = - 23'd255;
localparam signed [DEBIT:0]  W_2_x371 = - 23'd840;
localparam signed [DEBIT:0]  W_2_x372 = - 23'd771;
localparam signed [DEBIT:0]  W_2_x373 = - 23'd508;
localparam signed [DEBIT:0]  W_2_x374 = - 23'd416;
localparam signed [DEBIT:0]  W_2_x375 = - 23'd379;
localparam signed [DEBIT:0]  W_2_x376 = - 23'd401;
localparam signed [DEBIT:0]  W_2_x377 = - 23'd251;
localparam signed [DEBIT:0]  W_2_x378 = - 23'd301;
localparam signed [DEBIT:0]  W_2_x379 = - 23'd332;
localparam signed [DEBIT:0]  W_2_x380 = - 23'd309;
localparam signed [DEBIT:0]  W_2_x381 = - 23'd227;
localparam signed [DEBIT:0]  W_2_x382 = - 23'd192;
localparam signed [DEBIT:0]  W_2_x383 = - 23'd205;
localparam signed [DEBIT:0]  W_2_x384 = - 23'd158;
localparam signed [DEBIT:0]  W_2_x385 = - 23'd150;
localparam signed [DEBIT:0]  W_2_x386 = - 23'd349;
localparam signed [DEBIT:0]  W_2_x387 = - 23'd445;
localparam signed [DEBIT:0]  W_2_x388 = - 23'd267;
localparam signed [DEBIT:0]  W_2_x389 =  23'd333;
localparam signed [DEBIT:0]  W_2_x390 =  23'd894;
localparam signed [DEBIT:0]  W_2_x391 =  23'd974;
localparam signed [DEBIT:0]  W_2_x392 =  23'd982;
localparam signed [DEBIT:0]  W_2_x393 =  23'd971;
localparam signed [DEBIT:0]  W_2_x394 =  23'd952;
localparam signed [DEBIT:0]  W_2_x395 =  23'd949;
localparam signed [DEBIT:0]  W_2_x396 =  23'd795;
localparam signed [DEBIT:0]  W_2_x397 =  23'd506;
localparam signed [DEBIT:0]  W_2_x398 = - 23'd194;
localparam signed [DEBIT:0]  W_2_x399 = - 23'd632;
localparam signed [DEBIT:0]  W_2_x400 = - 23'd516;
localparam signed [DEBIT:0]  W_2_x401 = - 23'd311;
localparam signed [DEBIT:0]  W_2_x402 = - 23'd93;
localparam signed [DEBIT:0]  W_2_x403 = - 23'd45;
localparam signed [DEBIT:0]  W_2_x404 =  23'd18;
localparam signed [DEBIT:0]  W_2_x405 =  23'd60;
localparam signed [DEBIT:0]  W_2_x406 =  23'd44;
localparam signed [DEBIT:0]  W_2_x407 = - 23'd60;
localparam signed [DEBIT:0]  W_2_x408 = - 23'd230;
localparam signed [DEBIT:0]  W_2_x409 = - 23'd126;
localparam signed [DEBIT:0]  W_2_x410 = - 23'd295;
localparam signed [DEBIT:0]  W_2_x411 = - 23'd341;
localparam signed [DEBIT:0]  W_2_x412 = - 23'd261;
localparam signed [DEBIT:0]  W_2_x413 = - 23'd229;
localparam signed [DEBIT:0]  W_2_x414 = - 23'd363;
localparam signed [DEBIT:0]  W_2_x415 = - 23'd430;
localparam signed [DEBIT:0]  W_2_x416 = - 23'd342;
localparam signed [DEBIT:0]  W_2_x417 =  23'd237;
localparam signed [DEBIT:0]  W_2_x418 =  23'd834;
localparam signed [DEBIT:0]  W_2_x419 =  23'd979;
localparam signed [DEBIT:0]  W_2_x420 =  23'd962;
localparam signed [DEBIT:0]  W_2_x421 =  23'd972;
localparam signed [DEBIT:0]  W_2_x422 =  23'd960;
localparam signed [DEBIT:0]  W_2_x423 =  23'd942;
localparam signed [DEBIT:0]  W_2_x424 =  23'd826;
localparam signed [DEBIT:0]  W_2_x425 =  23'd572;
localparam signed [DEBIT:0]  W_2_x426 =  23'd63;
localparam signed [DEBIT:0]  W_2_x427 = - 23'd311;
localparam signed [DEBIT:0]  W_2_x428 = - 23'd235;
localparam signed [DEBIT:0]  W_2_x429 = - 23'd60;
localparam signed [DEBIT:0]  W_2_x430 =  23'd136;
localparam signed [DEBIT:0]  W_2_x431 =  23'd93;
localparam signed [DEBIT:0]  W_2_x432 =  23'd91;
localparam signed [DEBIT:0]  W_2_x433 =  23'd101;
localparam signed [DEBIT:0]  W_2_x434 =  23'd66;
localparam signed [DEBIT:0]  W_2_x435 = - 23'd97;
localparam signed [DEBIT:0]  W_2_x436 = - 23'd141;
localparam signed [DEBIT:0]  W_2_x437 = - 23'd103;
localparam signed [DEBIT:0]  W_2_x438 = - 23'd171;
localparam signed [DEBIT:0]  W_2_x439 = - 23'd252;
localparam signed [DEBIT:0]  W_2_x440 = - 23'd248;
localparam signed [DEBIT:0]  W_2_x441 = - 23'd348;
localparam signed [DEBIT:0]  W_2_x442 = - 23'd274;
localparam signed [DEBIT:0]  W_2_x443 = - 23'd360;
localparam signed [DEBIT:0]  W_2_x444 = - 23'd261;
localparam signed [DEBIT:0]  W_2_x445 =  23'd282;
localparam signed [DEBIT:0]  W_2_x446 =  23'd852;
localparam signed [DEBIT:0]  W_2_x447 =  23'd996;
localparam signed [DEBIT:0]  W_2_x448 =  23'd972;
localparam signed [DEBIT:0]  W_2_x449 =  23'd972;
localparam signed [DEBIT:0]  W_2_x450 =  23'd965;
localparam signed [DEBIT:0]  W_2_x451 =  23'd925;
localparam signed [DEBIT:0]  W_2_x452 =  23'd832;
localparam signed [DEBIT:0]  W_2_x453 =  23'd657;
localparam signed [DEBIT:0]  W_2_x454 =  23'd285;
localparam signed [DEBIT:0]  W_2_x455 =  23'd55;
localparam signed [DEBIT:0]  W_2_x456 = - 23'd10;
localparam signed [DEBIT:0]  W_2_x457 =  23'd54;
localparam signed [DEBIT:0]  W_2_x458 =  23'd98;
localparam signed [DEBIT:0]  W_2_x459 =  23'd111;
localparam signed [DEBIT:0]  W_2_x460 =  23'd179;
localparam signed [DEBIT:0]  W_2_x461 =  23'd229;
localparam signed [DEBIT:0]  W_2_x462 =  23'd179;
localparam signed [DEBIT:0]  W_2_x463 = - 23'd65;
localparam signed [DEBIT:0]  W_2_x464 =  23'd31;
localparam signed [DEBIT:0]  W_2_x465 =  23'd97;
localparam signed [DEBIT:0]  W_2_x466 =  23'd96;
localparam signed [DEBIT:0]  W_2_x467 = - 23'd57;
localparam signed [DEBIT:0]  W_2_x468 = - 23'd146;
localparam signed [DEBIT:0]  W_2_x469 = - 23'd151;
localparam signed [DEBIT:0]  W_2_x470 = - 23'd91;
localparam signed [DEBIT:0]  W_2_x471 = - 23'd112;
localparam signed [DEBIT:0]  W_2_x472 =  23'd2;
localparam signed [DEBIT:0]  W_2_x473 =  23'd450;
localparam signed [DEBIT:0]  W_2_x474 =  23'd974;
localparam signed [DEBIT:0]  W_2_x475 =  23'd1016;
localparam signed [DEBIT:0]  W_2_x476 =  23'd962;
localparam signed [DEBIT:0]  W_2_x477 =  23'd964;
localparam signed [DEBIT:0]  W_2_x478 =  23'd969;
localparam signed [DEBIT:0]  W_2_x479 =  23'd916;
localparam signed [DEBIT:0]  W_2_x480 =  23'd776;
localparam signed [DEBIT:0]  W_2_x481 =  23'd633;
localparam signed [DEBIT:0]  W_2_x482 =  23'd407;
localparam signed [DEBIT:0]  W_2_x483 =  23'd300;
localparam signed [DEBIT:0]  W_2_x484 =  23'd202;
localparam signed [DEBIT:0]  W_2_x485 =  23'd157;
localparam signed [DEBIT:0]  W_2_x486 =  23'd89;
localparam signed [DEBIT:0]  W_2_x487 =  23'd72;
localparam signed [DEBIT:0]  W_2_x488 =  23'd103;
localparam signed [DEBIT:0]  W_2_x489 =  23'd313;
localparam signed [DEBIT:0]  W_2_x490 =  23'd168;
localparam signed [DEBIT:0]  W_2_x491 =  23'd66;
localparam signed [DEBIT:0]  W_2_x492 =  23'd279;
localparam signed [DEBIT:0]  W_2_x493 =  23'd239;
localparam signed [DEBIT:0]  W_2_x494 =  23'd155;
localparam signed [DEBIT:0]  W_2_x495 = - 23'd70;
localparam signed [DEBIT:0]  W_2_x496 = - 23'd155;
localparam signed [DEBIT:0]  W_2_x497 = - 23'd96;
localparam signed [DEBIT:0]  W_2_x498 = - 23'd11;
localparam signed [DEBIT:0]  W_2_x499 =  23'd84;
localparam signed [DEBIT:0]  W_2_x500 =  23'd295;
localparam signed [DEBIT:0]  W_2_x501 =  23'd721;
localparam signed [DEBIT:0]  W_2_x502 =  23'd1044;
localparam signed [DEBIT:0]  W_2_x503 =  23'd1013;
localparam signed [DEBIT:0]  W_2_x504 =  23'd959;
localparam signed [DEBIT:0]  W_2_x505 =  23'd960;
localparam signed [DEBIT:0]  W_2_x506 =  23'd961;
localparam signed [DEBIT:0]  W_2_x507 =  23'd891;
localparam signed [DEBIT:0]  W_2_x508 =  23'd721;
localparam signed [DEBIT:0]  W_2_x509 =  23'd620;
localparam signed [DEBIT:0]  W_2_x510 =  23'd414;
localparam signed [DEBIT:0]  W_2_x511 =  23'd415;
localparam signed [DEBIT:0]  W_2_x512 =  23'd373;
localparam signed [DEBIT:0]  W_2_x513 =  23'd234;
localparam signed [DEBIT:0]  W_2_x514 =  23'd123;
localparam signed [DEBIT:0]  W_2_x515 =  23'd41;
localparam signed [DEBIT:0]  W_2_x516 =  23'd111;
localparam signed [DEBIT:0]  W_2_x517 =  23'd265;
localparam signed [DEBIT:0]  W_2_x518 =  23'd288;
localparam signed [DEBIT:0]  W_2_x519 =  23'd261;
localparam signed [DEBIT:0]  W_2_x520 =  23'd85;
localparam signed [DEBIT:0]  W_2_x521 =  23'd71;
localparam signed [DEBIT:0]  W_2_x522 = - 23'd24;
localparam signed [DEBIT:0]  W_2_x523 = - 23'd90;
localparam signed [DEBIT:0]  W_2_x524 = - 23'd183;
localparam signed [DEBIT:0]  W_2_x525 = - 23'd103;
localparam signed [DEBIT:0]  W_2_x526 =  23'd3;
localparam signed [DEBIT:0]  W_2_x527 =  23'd114;
localparam signed [DEBIT:0]  W_2_x528 =  23'd516;
localparam signed [DEBIT:0]  W_2_x529 =  23'd916;
localparam signed [DEBIT:0]  W_2_x530 =  23'd1030;
localparam signed [DEBIT:0]  W_2_x531 =  23'd976;
localparam signed [DEBIT:0]  W_2_x532 =  23'd972;
localparam signed [DEBIT:0]  W_2_x533 =  23'd970;
localparam signed [DEBIT:0]  W_2_x534 =  23'd959;
localparam signed [DEBIT:0]  W_2_x535 =  23'd890;
localparam signed [DEBIT:0]  W_2_x536 =  23'd639;
localparam signed [DEBIT:0]  W_2_x537 =  23'd542;
localparam signed [DEBIT:0]  W_2_x538 =  23'd377;
localparam signed [DEBIT:0]  W_2_x539 =  23'd354;
localparam signed [DEBIT:0]  W_2_x540 =  23'd318;
localparam signed [DEBIT:0]  W_2_x541 =  23'd254;
localparam signed [DEBIT:0]  W_2_x542 =  23'd249;
localparam signed [DEBIT:0]  W_2_x543 =  23'd169;
localparam signed [DEBIT:0]  W_2_x544 =  23'd152;
localparam signed [DEBIT:0]  W_2_x545 =  23'd142;
localparam signed [DEBIT:0]  W_2_x546 =  23'd130;
localparam signed [DEBIT:0]  W_2_x547 =  23'd122;
localparam signed [DEBIT:0]  W_2_x548 =  23'd80;
localparam signed [DEBIT:0]  W_2_x549 = - 23'd47;
localparam signed [DEBIT:0]  W_2_x550 = - 23'd99;
localparam signed [DEBIT:0]  W_2_x551 = - 23'd103;
localparam signed [DEBIT:0]  W_2_x552 = - 23'd83;
localparam signed [DEBIT:0]  W_2_x553 = - 23'd89;
localparam signed [DEBIT:0]  W_2_x554 = - 23'd54;
localparam signed [DEBIT:0]  W_2_x555 =  23'd151;
localparam signed [DEBIT:0]  W_2_x556 =  23'd655;
localparam signed [DEBIT:0]  W_2_x557 =  23'd991;
localparam signed [DEBIT:0]  W_2_x558 =  23'd1020;
localparam signed [DEBIT:0]  W_2_x559 =  23'd959;
localparam signed [DEBIT:0]  W_2_x560 =  23'd962;
localparam signed [DEBIT:0]  W_2_x561 =  23'd974;
localparam signed [DEBIT:0]  W_2_x562 =  23'd950;
localparam signed [DEBIT:0]  W_2_x563 =  23'd895;
localparam signed [DEBIT:0]  W_2_x564 =  23'd664;
localparam signed [DEBIT:0]  W_2_x565 =  23'd468;
localparam signed [DEBIT:0]  W_2_x566 =  23'd304;
localparam signed [DEBIT:0]  W_2_x567 =  23'd240;
localparam signed [DEBIT:0]  W_2_x568 =  23'd225;
localparam signed [DEBIT:0]  W_2_x569 =  23'd184;
localparam signed [DEBIT:0]  W_2_x570 =  23'd294;
localparam signed [DEBIT:0]  W_2_x571 =  23'd214;
localparam signed [DEBIT:0]  W_2_x572 =  23'd19;
localparam signed [DEBIT:0]  W_2_x573 = - 23'd249;
localparam signed [DEBIT:0]  W_2_x574 = - 23'd270;
localparam signed [DEBIT:0]  W_2_x575 = - 23'd219;
localparam signed [DEBIT:0]  W_2_x576 = - 23'd219;
localparam signed [DEBIT:0]  W_2_x577 = - 23'd98;
localparam signed [DEBIT:0]  W_2_x578 = - 23'd100;
localparam signed [DEBIT:0]  W_2_x579 = - 23'd25;
localparam signed [DEBIT:0]  W_2_x580 = - 23'd27;
localparam signed [DEBIT:0]  W_2_x581 = - 23'd112;
localparam signed [DEBIT:0]  W_2_x582 =  23'd1;
localparam signed [DEBIT:0]  W_2_x583 =  23'd284;
localparam signed [DEBIT:0]  W_2_x584 =  23'd765;
localparam signed [DEBIT:0]  W_2_x585 =  23'd986;
localparam signed [DEBIT:0]  W_2_x586 =  23'd1009;
localparam signed [DEBIT:0]  W_2_x587 =  23'd966;
localparam signed [DEBIT:0]  W_2_x588 =  23'd963;
localparam signed [DEBIT:0]  W_2_x589 =  23'd967;
localparam signed [DEBIT:0]  W_2_x590 =  23'd960;
localparam signed [DEBIT:0]  W_2_x591 =  23'd910;
localparam signed [DEBIT:0]  W_2_x592 =  23'd741;
localparam signed [DEBIT:0]  W_2_x593 =  23'd457;
localparam signed [DEBIT:0]  W_2_x594 =  23'd201;
localparam signed [DEBIT:0]  W_2_x595 =  23'd45;
localparam signed [DEBIT:0]  W_2_x596 =  23'd7;
localparam signed [DEBIT:0]  W_2_x597 =  23'd69;
localparam signed [DEBIT:0]  W_2_x598 =  23'd124;
localparam signed [DEBIT:0]  W_2_x599 =  23'd81;
localparam signed [DEBIT:0]  W_2_x600 =  23'd29;
localparam signed [DEBIT:0]  W_2_x601 = - 23'd156;
localparam signed [DEBIT:0]  W_2_x602 = - 23'd196;
localparam signed [DEBIT:0]  W_2_x603 = - 23'd194;
localparam signed [DEBIT:0]  W_2_x604 = - 23'd154;
localparam signed [DEBIT:0]  W_2_x605 = - 23'd66;
localparam signed [DEBIT:0]  W_2_x606 =  23'd45;
localparam signed [DEBIT:0]  W_2_x607 =  23'd146;
localparam signed [DEBIT:0]  W_2_x608 =  23'd86;
localparam signed [DEBIT:0]  W_2_x609 = - 23'd30;
localparam signed [DEBIT:0]  W_2_x610 =  23'd96;
localparam signed [DEBIT:0]  W_2_x611 =  23'd415;
localparam signed [DEBIT:0]  W_2_x612 =  23'd810;
localparam signed [DEBIT:0]  W_2_x613 =  23'd905;
localparam signed [DEBIT:0]  W_2_x614 =  23'd964;
localparam signed [DEBIT:0]  W_2_x615 =  23'd949;
localparam signed [DEBIT:0]  W_2_x616 =  23'd966;
localparam signed [DEBIT:0]  W_2_x617 =  23'd966;
localparam signed [DEBIT:0]  W_2_x618 =  23'd962;
localparam signed [DEBIT:0]  W_2_x619 =  23'd913;
localparam signed [DEBIT:0]  W_2_x620 =  23'd815;
localparam signed [DEBIT:0]  W_2_x621 =  23'd581;
localparam signed [DEBIT:0]  W_2_x622 =  23'd217;
localparam signed [DEBIT:0]  W_2_x623 =  23'd9;
localparam signed [DEBIT:0]  W_2_x624 = - 23'd36;
localparam signed [DEBIT:0]  W_2_x625 =  23'd23;
localparam signed [DEBIT:0]  W_2_x626 =  23'd138;
localparam signed [DEBIT:0]  W_2_x627 =  23'd98;
localparam signed [DEBIT:0]  W_2_x628 =  23'd95;
localparam signed [DEBIT:0]  W_2_x629 =  23'd111;
localparam signed [DEBIT:0]  W_2_x630 = - 23'd24;
localparam signed [DEBIT:0]  W_2_x631 = - 23'd64;
localparam signed [DEBIT:0]  W_2_x632 = - 23'd98;
localparam signed [DEBIT:0]  W_2_x633 = - 23'd110;
localparam signed [DEBIT:0]  W_2_x634 = - 23'd36;
localparam signed [DEBIT:0]  W_2_x635 =  23'd83;
localparam signed [DEBIT:0]  W_2_x636 = - 23'd11;
localparam signed [DEBIT:0]  W_2_x637 =  23'd43;
localparam signed [DEBIT:0]  W_2_x638 =  23'd298;
localparam signed [DEBIT:0]  W_2_x639 =  23'd566;
localparam signed [DEBIT:0]  W_2_x640 =  23'd765;
localparam signed [DEBIT:0]  W_2_x641 =  23'd919;
localparam signed [DEBIT:0]  W_2_x642 =  23'd979;
localparam signed [DEBIT:0]  W_2_x643 =  23'd959;
localparam signed [DEBIT:0]  W_2_x644 =  23'd967;
localparam signed [DEBIT:0]  W_2_x645 =  23'd958;
localparam signed [DEBIT:0]  W_2_x646 =  23'd969;
localparam signed [DEBIT:0]  W_2_x647 =  23'd954;
localparam signed [DEBIT:0]  W_2_x648 =  23'd888;
localparam signed [DEBIT:0]  W_2_x649 =  23'd690;
localparam signed [DEBIT:0]  W_2_x650 =  23'd404;
localparam signed [DEBIT:0]  W_2_x651 =  23'd179;
localparam signed [DEBIT:0]  W_2_x652 =  23'd19;
localparam signed [DEBIT:0]  W_2_x653 = - 23'd79;
localparam signed [DEBIT:0]  W_2_x654 = - 23'd150;
localparam signed [DEBIT:0]  W_2_x655 = - 23'd184;
localparam signed [DEBIT:0]  W_2_x656 = - 23'd162;
localparam signed [DEBIT:0]  W_2_x657 = - 23'd133;
localparam signed [DEBIT:0]  W_2_x658 = - 23'd266;
localparam signed [DEBIT:0]  W_2_x659 = - 23'd308;
localparam signed [DEBIT:0]  W_2_x660 = - 23'd276;
localparam signed [DEBIT:0]  W_2_x661 = - 23'd252;
localparam signed [DEBIT:0]  W_2_x662 = - 23'd217;
localparam signed [DEBIT:0]  W_2_x663 = - 23'd73;
localparam signed [DEBIT:0]  W_2_x664 =  23'd113;
localparam signed [DEBIT:0]  W_2_x665 =  23'd235;
localparam signed [DEBIT:0]  W_2_x666 =  23'd489;
localparam signed [DEBIT:0]  W_2_x667 =  23'd693;
localparam signed [DEBIT:0]  W_2_x668 =  23'd835;
localparam signed [DEBIT:0]  W_2_x669 =  23'd939;
localparam signed [DEBIT:0]  W_2_x670 =  23'd970;
localparam signed [DEBIT:0]  W_2_x671 =  23'd966;
localparam signed [DEBIT:0]  W_2_x672 =  23'd960;
localparam signed [DEBIT:0]  W_2_x673 =  23'd964;
localparam signed [DEBIT:0]  W_2_x674 =  23'd965;
localparam signed [DEBIT:0]  W_2_x675 =  23'd951;
localparam signed [DEBIT:0]  W_2_x676 =  23'd910;
localparam signed [DEBIT:0]  W_2_x677 =  23'd776;
localparam signed [DEBIT:0]  W_2_x678 =  23'd622;
localparam signed [DEBIT:0]  W_2_x679 =  23'd447;
localparam signed [DEBIT:0]  W_2_x680 =  23'd248;
localparam signed [DEBIT:0]  W_2_x681 =  23'd95;
localparam signed [DEBIT:0]  W_2_x682 = - 23'd88;
localparam signed [DEBIT:0]  W_2_x683 = - 23'd162;
localparam signed [DEBIT:0]  W_2_x684 = - 23'd66;
localparam signed [DEBIT:0]  W_2_x685 = - 23'd2;
localparam signed [DEBIT:0]  W_2_x686 =  23'd33;
localparam signed [DEBIT:0]  W_2_x687 =  23'd1;
localparam signed [DEBIT:0]  W_2_x688 = - 23'd63;
localparam signed [DEBIT:0]  W_2_x689 = - 23'd75;
localparam signed [DEBIT:0]  W_2_x690 =  23'd59;
localparam signed [DEBIT:0]  W_2_x691 =  23'd202;
localparam signed [DEBIT:0]  W_2_x692 =  23'd340;
localparam signed [DEBIT:0]  W_2_x693 =  23'd418;
localparam signed [DEBIT:0]  W_2_x694 =  23'd578;
localparam signed [DEBIT:0]  W_2_x695 =  23'd750;
localparam signed [DEBIT:0]  W_2_x696 =  23'd879;
localparam signed [DEBIT:0]  W_2_x697 =  23'd973;
localparam signed [DEBIT:0]  W_2_x698 =  23'd972;
localparam signed [DEBIT:0]  W_2_x699 =  23'd976;
localparam signed [DEBIT:0]  W_2_x700 =  23'd970;
localparam signed [DEBIT:0]  W_2_x701 =  23'd962;
localparam signed [DEBIT:0]  W_2_x702 =  23'd963;
localparam signed [DEBIT:0]  W_2_x703 =  23'd965;
localparam signed [DEBIT:0]  W_2_x704 =  23'd946;
localparam signed [DEBIT:0]  W_2_x705 =  23'd886;
localparam signed [DEBIT:0]  W_2_x706 =  23'd831;
localparam signed [DEBIT:0]  W_2_x707 =  23'd746;
localparam signed [DEBIT:0]  W_2_x708 =  23'd636;
localparam signed [DEBIT:0]  W_2_x709 =  23'd528;
localparam signed [DEBIT:0]  W_2_x710 =  23'd438;
localparam signed [DEBIT:0]  W_2_x711 =  23'd415;
localparam signed [DEBIT:0]  W_2_x712 =  23'd426;
localparam signed [DEBIT:0]  W_2_x713 =  23'd416;
localparam signed [DEBIT:0]  W_2_x714 =  23'd434;
localparam signed [DEBIT:0]  W_2_x715 =  23'd457;
localparam signed [DEBIT:0]  W_2_x716 =  23'd466;
localparam signed [DEBIT:0]  W_2_x717 =  23'd445;
localparam signed [DEBIT:0]  W_2_x718 =  23'd514;
localparam signed [DEBIT:0]  W_2_x719 =  23'd564;
localparam signed [DEBIT:0]  W_2_x720 =  23'd625;
localparam signed [DEBIT:0]  W_2_x721 =  23'd661;
localparam signed [DEBIT:0]  W_2_x722 =  23'd738;
localparam signed [DEBIT:0]  W_2_x723 =  23'd826;
localparam signed [DEBIT:0]  W_2_x724 =  23'd915;
localparam signed [DEBIT:0]  W_2_x725 =  23'd955;
localparam signed [DEBIT:0]  W_2_x726 =  23'd968;
localparam signed [DEBIT:0]  W_2_x727 =  23'd969;
localparam signed [DEBIT:0]  W_2_x728 =  23'd973;
localparam signed [DEBIT:0]  W_2_x729 =  23'd970;
localparam signed [DEBIT:0]  W_2_x730 =  23'd975;
localparam signed [DEBIT:0]  W_2_x731 =  23'd967;
localparam signed [DEBIT:0]  W_2_x732 =  23'd970;
localparam signed [DEBIT:0]  W_2_x733 =  23'd968;
localparam signed [DEBIT:0]  W_2_x734 =  23'd941;
localparam signed [DEBIT:0]  W_2_x735 =  23'd897;
localparam signed [DEBIT:0]  W_2_x736 =  23'd845;
localparam signed [DEBIT:0]  W_2_x737 =  23'd797;
localparam signed [DEBIT:0]  W_2_x738 =  23'd783;
localparam signed [DEBIT:0]  W_2_x739 =  23'd766;
localparam signed [DEBIT:0]  W_2_x740 =  23'd773;
localparam signed [DEBIT:0]  W_2_x741 =  23'd777;
localparam signed [DEBIT:0]  W_2_x742 =  23'd735;
localparam signed [DEBIT:0]  W_2_x743 =  23'd718;
localparam signed [DEBIT:0]  W_2_x744 =  23'd704;
localparam signed [DEBIT:0]  W_2_x745 =  23'd634;
localparam signed [DEBIT:0]  W_2_x746 =  23'd682;
localparam signed [DEBIT:0]  W_2_x747 =  23'd727;
localparam signed [DEBIT:0]  W_2_x748 =  23'd812;
localparam signed [DEBIT:0]  W_2_x749 =  23'd840;
localparam signed [DEBIT:0]  W_2_x750 =  23'd875;
localparam signed [DEBIT:0]  W_2_x751 =  23'd922;
localparam signed [DEBIT:0]  W_2_x752 =  23'd948;
localparam signed [DEBIT:0]  W_2_x753 =  23'd968;
localparam signed [DEBIT:0]  W_2_x754 =  23'd965;
localparam signed [DEBIT:0]  W_2_x755 =  23'd965;
localparam signed [DEBIT:0]  W_2_x756 =  23'd970;
localparam signed [DEBIT:0]  W_2_x757 =  23'd965;
localparam signed [DEBIT:0]  W_2_x758 =  23'd966;
localparam signed [DEBIT:0]  W_2_x759 =  23'd974;
localparam signed [DEBIT:0]  W_2_x760 =  23'd972;
localparam signed [DEBIT:0]  W_2_x761 =  23'd969;
localparam signed [DEBIT:0]  W_2_x762 =  23'd964;
localparam signed [DEBIT:0]  W_2_x763 =  23'd947;
localparam signed [DEBIT:0]  W_2_x764 =  23'd950;
localparam signed [DEBIT:0]  W_2_x765 =  23'd952;
localparam signed [DEBIT:0]  W_2_x766 =  23'd965;
localparam signed [DEBIT:0]  W_2_x767 =  23'd952;
localparam signed [DEBIT:0]  W_2_x768 =  23'd945;
localparam signed [DEBIT:0]  W_2_x769 =  23'd935;
localparam signed [DEBIT:0]  W_2_x770 =  23'd939;
localparam signed [DEBIT:0]  W_2_x771 =  23'd919;
localparam signed [DEBIT:0]  W_2_x772 =  23'd881;
localparam signed [DEBIT:0]  W_2_x773 =  23'd879;
localparam signed [DEBIT:0]  W_2_x774 =  23'd888;
localparam signed [DEBIT:0]  W_2_x775 =  23'd907;
localparam signed [DEBIT:0]  W_2_x776 =  23'd934;
localparam signed [DEBIT:0]  W_2_x777 =  23'd939;
localparam signed [DEBIT:0]  W_2_x778 =  23'd953;
localparam signed [DEBIT:0]  W_2_x779 =  23'd945;
localparam signed [DEBIT:0]  W_2_x780 =  23'd972;
localparam signed [DEBIT:0]  W_2_x781 =  23'd976;
localparam signed [DEBIT:0]  W_2_x782 =  23'd958;
localparam signed [DEBIT:0]  W_2_x783 =  23'd965;
localparam signed [DEBIT:0]  W_2_x784 =  23'd961;
localparam signed [DEBIT:0]  W_3_x1 =  23'd965;
localparam signed [DEBIT:0]  W_3_x2 =  23'd963;
localparam signed [DEBIT:0]  W_3_x3 =  23'd957;
localparam signed [DEBIT:0]  W_3_x4 =  23'd962;
localparam signed [DEBIT:0]  W_3_x5 =  23'd956;
localparam signed [DEBIT:0]  W_3_x6 =  23'd960;
localparam signed [DEBIT:0]  W_3_x7 =  23'd965;
localparam signed [DEBIT:0]  W_3_x8 =  23'd962;
localparam signed [DEBIT:0]  W_3_x9 =  23'd965;
localparam signed [DEBIT:0]  W_3_x10 =  23'd968;
localparam signed [DEBIT:0]  W_3_x11 =  23'd961;
localparam signed [DEBIT:0]  W_3_x12 =  23'd958;
localparam signed [DEBIT:0]  W_3_x13 =  23'd964;
localparam signed [DEBIT:0]  W_3_x14 =  23'd962;
localparam signed [DEBIT:0]  W_3_x15 =  23'd960;
localparam signed [DEBIT:0]  W_3_x16 =  23'd959;
localparam signed [DEBIT:0]  W_3_x17 =  23'd959;
localparam signed [DEBIT:0]  W_3_x18 =  23'd966;
localparam signed [DEBIT:0]  W_3_x19 =  23'd957;
localparam signed [DEBIT:0]  W_3_x20 =  23'd963;
localparam signed [DEBIT:0]  W_3_x21 =  23'd964;
localparam signed [DEBIT:0]  W_3_x22 =  23'd951;
localparam signed [DEBIT:0]  W_3_x23 =  23'd963;
localparam signed [DEBIT:0]  W_3_x24 =  23'd967;
localparam signed [DEBIT:0]  W_3_x25 =  23'd966;
localparam signed [DEBIT:0]  W_3_x26 =  23'd960;
localparam signed [DEBIT:0]  W_3_x27 =  23'd962;
localparam signed [DEBIT:0]  W_3_x28 =  23'd958;
localparam signed [DEBIT:0]  W_3_x29 =  23'd972;
localparam signed [DEBIT:0]  W_3_x30 =  23'd964;
localparam signed [DEBIT:0]  W_3_x31 =  23'd964;
localparam signed [DEBIT:0]  W_3_x32 =  23'd960;
localparam signed [DEBIT:0]  W_3_x33 =  23'd961;
localparam signed [DEBIT:0]  W_3_x34 =  23'd962;
localparam signed [DEBIT:0]  W_3_x35 =  23'd965;
localparam signed [DEBIT:0]  W_3_x36 =  23'd961;
localparam signed [DEBIT:0]  W_3_x37 =  23'd958;
localparam signed [DEBIT:0]  W_3_x38 =  23'd964;
localparam signed [DEBIT:0]  W_3_x39 =  23'd943;
localparam signed [DEBIT:0]  W_3_x40 =  23'd938;
localparam signed [DEBIT:0]  W_3_x41 =  23'd947;
localparam signed [DEBIT:0]  W_3_x42 =  23'd948;
localparam signed [DEBIT:0]  W_3_x43 =  23'd948;
localparam signed [DEBIT:0]  W_3_x44 =  23'd953;
localparam signed [DEBIT:0]  W_3_x45 =  23'd953;
localparam signed [DEBIT:0]  W_3_x46 =  23'd971;
localparam signed [DEBIT:0]  W_3_x47 =  23'd961;
localparam signed [DEBIT:0]  W_3_x48 =  23'd962;
localparam signed [DEBIT:0]  W_3_x49 =  23'd961;
localparam signed [DEBIT:0]  W_3_x50 =  23'd967;
localparam signed [DEBIT:0]  W_3_x51 =  23'd967;
localparam signed [DEBIT:0]  W_3_x52 =  23'd965;
localparam signed [DEBIT:0]  W_3_x53 =  23'd957;
localparam signed [DEBIT:0]  W_3_x54 =  23'd961;
localparam signed [DEBIT:0]  W_3_x55 =  23'd965;
localparam signed [DEBIT:0]  W_3_x56 =  23'd959;
localparam signed [DEBIT:0]  W_3_x57 =  23'd951;
localparam signed [DEBIT:0]  W_3_x58 =  23'd957;
localparam signed [DEBIT:0]  W_3_x59 =  23'd962;
localparam signed [DEBIT:0]  W_3_x60 =  23'd966;
localparam signed [DEBIT:0]  W_3_x61 =  23'd961;
localparam signed [DEBIT:0]  W_3_x62 =  23'd961;
localparam signed [DEBIT:0]  W_3_x63 =  23'd963;
localparam signed [DEBIT:0]  W_3_x64 =  23'd941;
localparam signed [DEBIT:0]  W_3_x65 =  23'd922;
localparam signed [DEBIT:0]  W_3_x66 =  23'd872;
localparam signed [DEBIT:0]  W_3_x67 =  23'd860;
localparam signed [DEBIT:0]  W_3_x68 =  23'd847;
localparam signed [DEBIT:0]  W_3_x69 =  23'd828;
localparam signed [DEBIT:0]  W_3_x70 =  23'd815;
localparam signed [DEBIT:0]  W_3_x71 =  23'd800;
localparam signed [DEBIT:0]  W_3_x72 =  23'd829;
localparam signed [DEBIT:0]  W_3_x73 =  23'd840;
localparam signed [DEBIT:0]  W_3_x74 =  23'd871;
localparam signed [DEBIT:0]  W_3_x75 =  23'd898;
localparam signed [DEBIT:0]  W_3_x76 =  23'd913;
localparam signed [DEBIT:0]  W_3_x77 =  23'd952;
localparam signed [DEBIT:0]  W_3_x78 =  23'd950;
localparam signed [DEBIT:0]  W_3_x79 =  23'd952;
localparam signed [DEBIT:0]  W_3_x80 =  23'd955;
localparam signed [DEBIT:0]  W_3_x81 =  23'd961;
localparam signed [DEBIT:0]  W_3_x82 =  23'd954;
localparam signed [DEBIT:0]  W_3_x83 =  23'd966;
localparam signed [DEBIT:0]  W_3_x84 =  23'd968;
localparam signed [DEBIT:0]  W_3_x85 =  23'd965;
localparam signed [DEBIT:0]  W_3_x86 =  23'd962;
localparam signed [DEBIT:0]  W_3_x87 =  23'd960;
localparam signed [DEBIT:0]  W_3_x88 =  23'd969;
localparam signed [DEBIT:0]  W_3_x89 =  23'd960;
localparam signed [DEBIT:0]  W_3_x90 =  23'd958;
localparam signed [DEBIT:0]  W_3_x91 =  23'd910;
localparam signed [DEBIT:0]  W_3_x92 =  23'd788;
localparam signed [DEBIT:0]  W_3_x93 =  23'd634;
localparam signed [DEBIT:0]  W_3_x94 =  23'd521;
localparam signed [DEBIT:0]  W_3_x95 =  23'd401;
localparam signed [DEBIT:0]  W_3_x96 =  23'd315;
localparam signed [DEBIT:0]  W_3_x97 =  23'd320;
localparam signed [DEBIT:0]  W_3_x98 =  23'd357;
localparam signed [DEBIT:0]  W_3_x99 =  23'd383;
localparam signed [DEBIT:0]  W_3_x100 =  23'd362;
localparam signed [DEBIT:0]  W_3_x101 =  23'd438;
localparam signed [DEBIT:0]  W_3_x102 =  23'd562;
localparam signed [DEBIT:0]  W_3_x103 =  23'd578;
localparam signed [DEBIT:0]  W_3_x104 =  23'd653;
localparam signed [DEBIT:0]  W_3_x105 =  23'd758;
localparam signed [DEBIT:0]  W_3_x106 =  23'd810;
localparam signed [DEBIT:0]  W_3_x107 =  23'd866;
localparam signed [DEBIT:0]  W_3_x108 =  23'd935;
localparam signed [DEBIT:0]  W_3_x109 =  23'd960;
localparam signed [DEBIT:0]  W_3_x110 =  23'd971;
localparam signed [DEBIT:0]  W_3_x111 =  23'd961;
localparam signed [DEBIT:0]  W_3_x112 =  23'd961;
localparam signed [DEBIT:0]  W_3_x113 =  23'd961;
localparam signed [DEBIT:0]  W_3_x114 =  23'd954;
localparam signed [DEBIT:0]  W_3_x115 =  23'd958;
localparam signed [DEBIT:0]  W_3_x116 =  23'd956;
localparam signed [DEBIT:0]  W_3_x117 =  23'd966;
localparam signed [DEBIT:0]  W_3_x118 =  23'd907;
localparam signed [DEBIT:0]  W_3_x119 =  23'd739;
localparam signed [DEBIT:0]  W_3_x120 =  23'd559;
localparam signed [DEBIT:0]  W_3_x121 =  23'd363;
localparam signed [DEBIT:0]  W_3_x122 =  23'd181;
localparam signed [DEBIT:0]  W_3_x123 =  23'd204;
localparam signed [DEBIT:0]  W_3_x124 =  23'd179;
localparam signed [DEBIT:0]  W_3_x125 =  23'd144;
localparam signed [DEBIT:0]  W_3_x126 =  23'd160;
localparam signed [DEBIT:0]  W_3_x127 =  23'd212;
localparam signed [DEBIT:0]  W_3_x128 =  23'd250;
localparam signed [DEBIT:0]  W_3_x129 =  23'd114;
localparam signed [DEBIT:0]  W_3_x130 =  23'd98;
localparam signed [DEBIT:0]  W_3_x131 =  23'd158;
localparam signed [DEBIT:0]  W_3_x132 =  23'd189;
localparam signed [DEBIT:0]  W_3_x133 =  23'd192;
localparam signed [DEBIT:0]  W_3_x134 =  23'd297;
localparam signed [DEBIT:0]  W_3_x135 =  23'd487;
localparam signed [DEBIT:0]  W_3_x136 =  23'd692;
localparam signed [DEBIT:0]  W_3_x137 =  23'd855;
localparam signed [DEBIT:0]  W_3_x138 =  23'd944;
localparam signed [DEBIT:0]  W_3_x139 =  23'd968;
localparam signed [DEBIT:0]  W_3_x140 =  23'd959;
localparam signed [DEBIT:0]  W_3_x141 =  23'd969;
localparam signed [DEBIT:0]  W_3_x142 =  23'd961;
localparam signed [DEBIT:0]  W_3_x143 =  23'd966;
localparam signed [DEBIT:0]  W_3_x144 =  23'd965;
localparam signed [DEBIT:0]  W_3_x145 =  23'd915;
localparam signed [DEBIT:0]  W_3_x146 =  23'd731;
localparam signed [DEBIT:0]  W_3_x147 =  23'd461;
localparam signed [DEBIT:0]  W_3_x148 =  23'd262;
localparam signed [DEBIT:0]  W_3_x149 =  23'd42;
localparam signed [DEBIT:0]  W_3_x150 =  23'd47;
localparam signed [DEBIT:0]  W_3_x151 =  23'd127;
localparam signed [DEBIT:0]  W_3_x152 =  23'd120;
localparam signed [DEBIT:0]  W_3_x153 =  23'd106;
localparam signed [DEBIT:0]  W_3_x154 =  23'd49;
localparam signed [DEBIT:0]  W_3_x155 =  23'd62;
localparam signed [DEBIT:0]  W_3_x156 =  23'd44;
localparam signed [DEBIT:0]  W_3_x157 =  23'd31;
localparam signed [DEBIT:0]  W_3_x158 = - 23'd181;
localparam signed [DEBIT:0]  W_3_x159 = - 23'd202;
localparam signed [DEBIT:0]  W_3_x160 = - 23'd231;
localparam signed [DEBIT:0]  W_3_x161 = - 23'd337;
localparam signed [DEBIT:0]  W_3_x162 = - 23'd343;
localparam signed [DEBIT:0]  W_3_x163 = - 23'd64;
localparam signed [DEBIT:0]  W_3_x164 =  23'd325;
localparam signed [DEBIT:0]  W_3_x165 =  23'd674;
localparam signed [DEBIT:0]  W_3_x166 =  23'd886;
localparam signed [DEBIT:0]  W_3_x167 =  23'd971;
localparam signed [DEBIT:0]  W_3_x168 =  23'd958;
localparam signed [DEBIT:0]  W_3_x169 =  23'd958;
localparam signed [DEBIT:0]  W_3_x170 =  23'd960;
localparam signed [DEBIT:0]  W_3_x171 =  23'd946;
localparam signed [DEBIT:0]  W_3_x172 =  23'd933;
localparam signed [DEBIT:0]  W_3_x173 =  23'd810;
localparam signed [DEBIT:0]  W_3_x174 =  23'd600;
localparam signed [DEBIT:0]  W_3_x175 =  23'd324;
localparam signed [DEBIT:0]  W_3_x176 =  23'd141;
localparam signed [DEBIT:0]  W_3_x177 =  23'd152;
localparam signed [DEBIT:0]  W_3_x178 =  23'd138;
localparam signed [DEBIT:0]  W_3_x179 =  23'd138;
localparam signed [DEBIT:0]  W_3_x180 =  23'd198;
localparam signed [DEBIT:0]  W_3_x181 =  23'd239;
localparam signed [DEBIT:0]  W_3_x182 =  23'd228;
localparam signed [DEBIT:0]  W_3_x183 =  23'd184;
localparam signed [DEBIT:0]  W_3_x184 =  23'd130;
localparam signed [DEBIT:0]  W_3_x185 =  23'd122;
localparam signed [DEBIT:0]  W_3_x186 =  23'd75;
localparam signed [DEBIT:0]  W_3_x187 = - 23'd13;
localparam signed [DEBIT:0]  W_3_x188 = - 23'd177;
localparam signed [DEBIT:0]  W_3_x189 = - 23'd266;
localparam signed [DEBIT:0]  W_3_x190 = - 23'd499;
localparam signed [DEBIT:0]  W_3_x191 = - 23'd345;
localparam signed [DEBIT:0]  W_3_x192 =  23'd84;
localparam signed [DEBIT:0]  W_3_x193 =  23'd488;
localparam signed [DEBIT:0]  W_3_x194 =  23'd793;
localparam signed [DEBIT:0]  W_3_x195 =  23'd934;
localparam signed [DEBIT:0]  W_3_x196 =  23'd957;
localparam signed [DEBIT:0]  W_3_x197 =  23'd954;
localparam signed [DEBIT:0]  W_3_x198 =  23'd967;
localparam signed [DEBIT:0]  W_3_x199 =  23'd883;
localparam signed [DEBIT:0]  W_3_x200 =  23'd779;
localparam signed [DEBIT:0]  W_3_x201 =  23'd615;
localparam signed [DEBIT:0]  W_3_x202 =  23'd305;
localparam signed [DEBIT:0]  W_3_x203 =  23'd63;
localparam signed [DEBIT:0]  W_3_x204 =  23'd23;
localparam signed [DEBIT:0]  W_3_x205 =  23'd75;
localparam signed [DEBIT:0]  W_3_x206 =  23'd74;
localparam signed [DEBIT:0]  W_3_x207 =  23'd79;
localparam signed [DEBIT:0]  W_3_x208 =  23'd83;
localparam signed [DEBIT:0]  W_3_x209 =  23'd143;
localparam signed [DEBIT:0]  W_3_x210 =  23'd107;
localparam signed [DEBIT:0]  W_3_x211 =  23'd102;
localparam signed [DEBIT:0]  W_3_x212 =  23'd144;
localparam signed [DEBIT:0]  W_3_x213 =  23'd35;
localparam signed [DEBIT:0]  W_3_x214 =  23'd81;
localparam signed [DEBIT:0]  W_3_x215 =  23'd115;
localparam signed [DEBIT:0]  W_3_x216 =  23'd124;
localparam signed [DEBIT:0]  W_3_x217 =  23'd11;
localparam signed [DEBIT:0]  W_3_x218 = - 23'd297;
localparam signed [DEBIT:0]  W_3_x219 = - 23'd305;
localparam signed [DEBIT:0]  W_3_x220 = - 23'd46;
localparam signed [DEBIT:0]  W_3_x221 =  23'd387;
localparam signed [DEBIT:0]  W_3_x222 =  23'd718;
localparam signed [DEBIT:0]  W_3_x223 =  23'd915;
localparam signed [DEBIT:0]  W_3_x224 =  23'd968;
localparam signed [DEBIT:0]  W_3_x225 =  23'd961;
localparam signed [DEBIT:0]  W_3_x226 =  23'd888;
localparam signed [DEBIT:0]  W_3_x227 =  23'd721;
localparam signed [DEBIT:0]  W_3_x228 =  23'd532;
localparam signed [DEBIT:0]  W_3_x229 =  23'd252;
localparam signed [DEBIT:0]  W_3_x230 = - 23'd9;
localparam signed [DEBIT:0]  W_3_x231 = - 23'd142;
localparam signed [DEBIT:0]  W_3_x232 = - 23'd74;
localparam signed [DEBIT:0]  W_3_x233 = - 23'd144;
localparam signed [DEBIT:0]  W_3_x234 = - 23'd69;
localparam signed [DEBIT:0]  W_3_x235 = - 23'd61;
localparam signed [DEBIT:0]  W_3_x236 = - 23'd81;
localparam signed [DEBIT:0]  W_3_x237 = - 23'd60;
localparam signed [DEBIT:0]  W_3_x238 = - 23'd181;
localparam signed [DEBIT:0]  W_3_x239 = - 23'd220;
localparam signed [DEBIT:0]  W_3_x240 = - 23'd136;
localparam signed [DEBIT:0]  W_3_x241 = - 23'd55;
localparam signed [DEBIT:0]  W_3_x242 = - 23'd3;
localparam signed [DEBIT:0]  W_3_x243 =  23'd68;
localparam signed [DEBIT:0]  W_3_x244 =  23'd198;
localparam signed [DEBIT:0]  W_3_x245 =  23'd113;
localparam signed [DEBIT:0]  W_3_x246 = - 23'd166;
localparam signed [DEBIT:0]  W_3_x247 = - 23'd209;
localparam signed [DEBIT:0]  W_3_x248 = - 23'd8;
localparam signed [DEBIT:0]  W_3_x249 =  23'd394;
localparam signed [DEBIT:0]  W_3_x250 =  23'd697;
localparam signed [DEBIT:0]  W_3_x251 =  23'd936;
localparam signed [DEBIT:0]  W_3_x252 =  23'd969;
localparam signed [DEBIT:0]  W_3_x253 =  23'd957;
localparam signed [DEBIT:0]  W_3_x254 =  23'd848;
localparam signed [DEBIT:0]  W_3_x255 =  23'd666;
localparam signed [DEBIT:0]  W_3_x256 =  23'd441;
localparam signed [DEBIT:0]  W_3_x257 =  23'd172;
localparam signed [DEBIT:0]  W_3_x258 = - 23'd142;
localparam signed [DEBIT:0]  W_3_x259 = - 23'd304;
localparam signed [DEBIT:0]  W_3_x260 = - 23'd225;
localparam signed [DEBIT:0]  W_3_x261 = - 23'd241;
localparam signed [DEBIT:0]  W_3_x262 = - 23'd239;
localparam signed [DEBIT:0]  W_3_x263 = - 23'd308;
localparam signed [DEBIT:0]  W_3_x264 = - 23'd442;
localparam signed [DEBIT:0]  W_3_x265 = - 23'd355;
localparam signed [DEBIT:0]  W_3_x266 = - 23'd212;
localparam signed [DEBIT:0]  W_3_x267 = - 23'd210;
localparam signed [DEBIT:0]  W_3_x268 = - 23'd80;
localparam signed [DEBIT:0]  W_3_x269 = - 23'd31;
localparam signed [DEBIT:0]  W_3_x270 = - 23'd36;
localparam signed [DEBIT:0]  W_3_x271 = - 23'd55;
localparam signed [DEBIT:0]  W_3_x272 =  23'd53;
localparam signed [DEBIT:0]  W_3_x273 =  23'd142;
localparam signed [DEBIT:0]  W_3_x274 = - 23'd170;
localparam signed [DEBIT:0]  W_3_x275 = - 23'd158;
localparam signed [DEBIT:0]  W_3_x276 =  23'd60;
localparam signed [DEBIT:0]  W_3_x277 =  23'd500;
localparam signed [DEBIT:0]  W_3_x278 =  23'd799;
localparam signed [DEBIT:0]  W_3_x279 =  23'd942;
localparam signed [DEBIT:0]  W_3_x280 =  23'd967;
localparam signed [DEBIT:0]  W_3_x281 =  23'd964;
localparam signed [DEBIT:0]  W_3_x282 =  23'd862;
localparam signed [DEBIT:0]  W_3_x283 =  23'd709;
localparam signed [DEBIT:0]  W_3_x284 =  23'd528;
localparam signed [DEBIT:0]  W_3_x285 =  23'd260;
localparam signed [DEBIT:0]  W_3_x286 = - 23'd70;
localparam signed [DEBIT:0]  W_3_x287 = - 23'd370;
localparam signed [DEBIT:0]  W_3_x288 = - 23'd389;
localparam signed [DEBIT:0]  W_3_x289 = - 23'd426;
localparam signed [DEBIT:0]  W_3_x290 = - 23'd441;
localparam signed [DEBIT:0]  W_3_x291 = - 23'd629;
localparam signed [DEBIT:0]  W_3_x292 = - 23'd636;
localparam signed [DEBIT:0]  W_3_x293 = - 23'd296;
localparam signed [DEBIT:0]  W_3_x294 = - 23'd12;
localparam signed [DEBIT:0]  W_3_x295 =  23'd169;
localparam signed [DEBIT:0]  W_3_x296 =  23'd212;
localparam signed [DEBIT:0]  W_3_x297 =  23'd94;
localparam signed [DEBIT:0]  W_3_x298 =  23'd20;
localparam signed [DEBIT:0]  W_3_x299 =  23'd2;
localparam signed [DEBIT:0]  W_3_x300 = - 23'd5;
localparam signed [DEBIT:0]  W_3_x301 =  23'd13;
localparam signed [DEBIT:0]  W_3_x302 = - 23'd93;
localparam signed [DEBIT:0]  W_3_x303 = - 23'd114;
localparam signed [DEBIT:0]  W_3_x304 =  23'd154;
localparam signed [DEBIT:0]  W_3_x305 =  23'd635;
localparam signed [DEBIT:0]  W_3_x306 =  23'd908;
localparam signed [DEBIT:0]  W_3_x307 =  23'd951;
localparam signed [DEBIT:0]  W_3_x308 =  23'd956;
localparam signed [DEBIT:0]  W_3_x309 =  23'd959;
localparam signed [DEBIT:0]  W_3_x310 =  23'd898;
localparam signed [DEBIT:0]  W_3_x311 =  23'd777;
localparam signed [DEBIT:0]  W_3_x312 =  23'd605;
localparam signed [DEBIT:0]  W_3_x313 =  23'd315;
localparam signed [DEBIT:0]  W_3_x314 = - 23'd100;
localparam signed [DEBIT:0]  W_3_x315 = - 23'd493;
localparam signed [DEBIT:0]  W_3_x316 = - 23'd553;
localparam signed [DEBIT:0]  W_3_x317 = - 23'd471;
localparam signed [DEBIT:0]  W_3_x318 = - 23'd419;
localparam signed [DEBIT:0]  W_3_x319 = - 23'd456;
localparam signed [DEBIT:0]  W_3_x320 = - 23'd327;
localparam signed [DEBIT:0]  W_3_x321 = - 23'd48;
localparam signed [DEBIT:0]  W_3_x322 =  23'd161;
localparam signed [DEBIT:0]  W_3_x323 =  23'd352;
localparam signed [DEBIT:0]  W_3_x324 =  23'd381;
localparam signed [DEBIT:0]  W_3_x325 =  23'd225;
localparam signed [DEBIT:0]  W_3_x326 =  23'd165;
localparam signed [DEBIT:0]  W_3_x327 =  23'd150;
localparam signed [DEBIT:0]  W_3_x328 =  23'd32;
localparam signed [DEBIT:0]  W_3_x329 = - 23'd102;
localparam signed [DEBIT:0]  W_3_x330 = - 23'd244;
localparam signed [DEBIT:0]  W_3_x331 = - 23'd199;
localparam signed [DEBIT:0]  W_3_x332 =  23'd149;
localparam signed [DEBIT:0]  W_3_x333 =  23'd640;
localparam signed [DEBIT:0]  W_3_x334 =  23'd915;
localparam signed [DEBIT:0]  W_3_x335 =  23'd946;
localparam signed [DEBIT:0]  W_3_x336 =  23'd972;
localparam signed [DEBIT:0]  W_3_x337 =  23'd955;
localparam signed [DEBIT:0]  W_3_x338 =  23'd925;
localparam signed [DEBIT:0]  W_3_x339 =  23'd847;
localparam signed [DEBIT:0]  W_3_x340 =  23'd693;
localparam signed [DEBIT:0]  W_3_x341 =  23'd379;
localparam signed [DEBIT:0]  W_3_x342 = - 23'd94;
localparam signed [DEBIT:0]  W_3_x343 = - 23'd494;
localparam signed [DEBIT:0]  W_3_x344 = - 23'd489;
localparam signed [DEBIT:0]  W_3_x345 = - 23'd244;
localparam signed [DEBIT:0]  W_3_x346 = - 23'd173;
localparam signed [DEBIT:0]  W_3_x347 = - 23'd220;
localparam signed [DEBIT:0]  W_3_x348 = - 23'd204;
localparam signed [DEBIT:0]  W_3_x349 =  23'd165;
localparam signed [DEBIT:0]  W_3_x350 =  23'd275;
localparam signed [DEBIT:0]  W_3_x351 =  23'd200;
localparam signed [DEBIT:0]  W_3_x352 =  23'd166;
localparam signed [DEBIT:0]  W_3_x353 =  23'd171;
localparam signed [DEBIT:0]  W_3_x354 =  23'd68;
localparam signed [DEBIT:0]  W_3_x355 =  23'd3;
localparam signed [DEBIT:0]  W_3_x356 = - 23'd103;
localparam signed [DEBIT:0]  W_3_x357 = - 23'd291;
localparam signed [DEBIT:0]  W_3_x358 = - 23'd309;
localparam signed [DEBIT:0]  W_3_x359 = - 23'd226;
localparam signed [DEBIT:0]  W_3_x360 =  23'd96;
localparam signed [DEBIT:0]  W_3_x361 =  23'd610;
localparam signed [DEBIT:0]  W_3_x362 =  23'd935;
localparam signed [DEBIT:0]  W_3_x363 =  23'd955;
localparam signed [DEBIT:0]  W_3_x364 =  23'd960;
localparam signed [DEBIT:0]  W_3_x365 =  23'd950;
localparam signed [DEBIT:0]  W_3_x366 =  23'd946;
localparam signed [DEBIT:0]  W_3_x367 =  23'd907;
localparam signed [DEBIT:0]  W_3_x368 =  23'd783;
localparam signed [DEBIT:0]  W_3_x369 =  23'd456;
localparam signed [DEBIT:0]  W_3_x370 = - 23'd23;
localparam signed [DEBIT:0]  W_3_x371 = - 23'd425;
localparam signed [DEBIT:0]  W_3_x372 = - 23'd408;
localparam signed [DEBIT:0]  W_3_x373 = - 23'd104;
localparam signed [DEBIT:0]  W_3_x374 = - 23'd53;
localparam signed [DEBIT:0]  W_3_x375 = - 23'd91;
localparam signed [DEBIT:0]  W_3_x376 = - 23'd17;
localparam signed [DEBIT:0]  W_3_x377 =  23'd293;
localparam signed [DEBIT:0]  W_3_x378 =  23'd163;
localparam signed [DEBIT:0]  W_3_x379 =  23'd15;
localparam signed [DEBIT:0]  W_3_x380 =  23'd42;
localparam signed [DEBIT:0]  W_3_x381 =  23'd259;
localparam signed [DEBIT:0]  W_3_x382 =  23'd91;
localparam signed [DEBIT:0]  W_3_x383 = - 23'd77;
localparam signed [DEBIT:0]  W_3_x384 = - 23'd122;
localparam signed [DEBIT:0]  W_3_x385 = - 23'd226;
localparam signed [DEBIT:0]  W_3_x386 = - 23'd233;
localparam signed [DEBIT:0]  W_3_x387 = - 23'd181;
localparam signed [DEBIT:0]  W_3_x388 =  23'd70;
localparam signed [DEBIT:0]  W_3_x389 =  23'd576;
localparam signed [DEBIT:0]  W_3_x390 =  23'd888;
localparam signed [DEBIT:0]  W_3_x391 =  23'd942;
localparam signed [DEBIT:0]  W_3_x392 =  23'd957;
localparam signed [DEBIT:0]  W_3_x393 =  23'd964;
localparam signed [DEBIT:0]  W_3_x394 =  23'd955;
localparam signed [DEBIT:0]  W_3_x395 =  23'd937;
localparam signed [DEBIT:0]  W_3_x396 =  23'd863;
localparam signed [DEBIT:0]  W_3_x397 =  23'd569;
localparam signed [DEBIT:0]  W_3_x398 =  23'd57;
localparam signed [DEBIT:0]  W_3_x399 = - 23'd346;
localparam signed [DEBIT:0]  W_3_x400 = - 23'd359;
localparam signed [DEBIT:0]  W_3_x401 = - 23'd108;
localparam signed [DEBIT:0]  W_3_x402 =  23'd16;
localparam signed [DEBIT:0]  W_3_x403 = - 23'd173;
localparam signed [DEBIT:0]  W_3_x404 = - 23'd17;
localparam signed [DEBIT:0]  W_3_x405 =  23'd145;
localparam signed [DEBIT:0]  W_3_x406 = - 23'd32;
localparam signed [DEBIT:0]  W_3_x407 = - 23'd29;
localparam signed [DEBIT:0]  W_3_x408 =  23'd117;
localparam signed [DEBIT:0]  W_3_x409 =  23'd173;
localparam signed [DEBIT:0]  W_3_x410 =  23'd17;
localparam signed [DEBIT:0]  W_3_x411 =  23'd0;
localparam signed [DEBIT:0]  W_3_x412 = - 23'd74;
localparam signed [DEBIT:0]  W_3_x413 = - 23'd14;
localparam signed [DEBIT:0]  W_3_x414 =  23'd25;
localparam signed [DEBIT:0]  W_3_x415 = - 23'd32;
localparam signed [DEBIT:0]  W_3_x416 =  23'd104;
localparam signed [DEBIT:0]  W_3_x417 =  23'd561;
localparam signed [DEBIT:0]  W_3_x418 =  23'd862;
localparam signed [DEBIT:0]  W_3_x419 =  23'd918;
localparam signed [DEBIT:0]  W_3_x420 =  23'd966;
localparam signed [DEBIT:0]  W_3_x421 =  23'd963;
localparam signed [DEBIT:0]  W_3_x422 =  23'd969;
localparam signed [DEBIT:0]  W_3_x423 =  23'd958;
localparam signed [DEBIT:0]  W_3_x424 =  23'd885;
localparam signed [DEBIT:0]  W_3_x425 =  23'd656;
localparam signed [DEBIT:0]  W_3_x426 =  23'd134;
localparam signed [DEBIT:0]  W_3_x427 = - 23'd269;
localparam signed [DEBIT:0]  W_3_x428 = - 23'd333;
localparam signed [DEBIT:0]  W_3_x429 = - 23'd229;
localparam signed [DEBIT:0]  W_3_x430 = - 23'd102;
localparam signed [DEBIT:0]  W_3_x431 = - 23'd137;
localparam signed [DEBIT:0]  W_3_x432 =  23'd75;
localparam signed [DEBIT:0]  W_3_x433 =  23'd221;
localparam signed [DEBIT:0]  W_3_x434 =  23'd124;
localparam signed [DEBIT:0]  W_3_x435 =  23'd84;
localparam signed [DEBIT:0]  W_3_x436 =  23'd43;
localparam signed [DEBIT:0]  W_3_x437 = - 23'd14;
localparam signed [DEBIT:0]  W_3_x438 = - 23'd92;
localparam signed [DEBIT:0]  W_3_x439 = - 23'd4;
localparam signed [DEBIT:0]  W_3_x440 =  23'd90;
localparam signed [DEBIT:0]  W_3_x441 =  23'd189;
localparam signed [DEBIT:0]  W_3_x442 =  23'd238;
localparam signed [DEBIT:0]  W_3_x443 =  23'd136;
localparam signed [DEBIT:0]  W_3_x444 =  23'd118;
localparam signed [DEBIT:0]  W_3_x445 =  23'd521;
localparam signed [DEBIT:0]  W_3_x446 =  23'd828;
localparam signed [DEBIT:0]  W_3_x447 =  23'd917;
localparam signed [DEBIT:0]  W_3_x448 =  23'd959;
localparam signed [DEBIT:0]  W_3_x449 =  23'd964;
localparam signed [DEBIT:0]  W_3_x450 =  23'd955;
localparam signed [DEBIT:0]  W_3_x451 =  23'd978;
localparam signed [DEBIT:0]  W_3_x452 =  23'd938;
localparam signed [DEBIT:0]  W_3_x453 =  23'd689;
localparam signed [DEBIT:0]  W_3_x454 =  23'd120;
localparam signed [DEBIT:0]  W_3_x455 = - 23'd258;
localparam signed [DEBIT:0]  W_3_x456 = - 23'd297;
localparam signed [DEBIT:0]  W_3_x457 = - 23'd248;
localparam signed [DEBIT:0]  W_3_x458 = - 23'd217;
localparam signed [DEBIT:0]  W_3_x459 = - 23'd230;
localparam signed [DEBIT:0]  W_3_x460 = - 23'd111;
localparam signed [DEBIT:0]  W_3_x461 = - 23'd8;
localparam signed [DEBIT:0]  W_3_x462 = - 23'd60;
localparam signed [DEBIT:0]  W_3_x463 = - 23'd198;
localparam signed [DEBIT:0]  W_3_x464 = - 23'd135;
localparam signed [DEBIT:0]  W_3_x465 = - 23'd130;
localparam signed [DEBIT:0]  W_3_x466 = - 23'd6;
localparam signed [DEBIT:0]  W_3_x467 =  23'd43;
localparam signed [DEBIT:0]  W_3_x468 =  23'd116;
localparam signed [DEBIT:0]  W_3_x469 =  23'd247;
localparam signed [DEBIT:0]  W_3_x470 =  23'd228;
localparam signed [DEBIT:0]  W_3_x471 =  23'd217;
localparam signed [DEBIT:0]  W_3_x472 =  23'd172;
localparam signed [DEBIT:0]  W_3_x473 =  23'd433;
localparam signed [DEBIT:0]  W_3_x474 =  23'd758;
localparam signed [DEBIT:0]  W_3_x475 =  23'd920;
localparam signed [DEBIT:0]  W_3_x476 =  23'd955;
localparam signed [DEBIT:0]  W_3_x477 =  23'd958;
localparam signed [DEBIT:0]  W_3_x478 =  23'd960;
localparam signed [DEBIT:0]  W_3_x479 =  23'd983;
localparam signed [DEBIT:0]  W_3_x480 =  23'd990;
localparam signed [DEBIT:0]  W_3_x481 =  23'd698;
localparam signed [DEBIT:0]  W_3_x482 =  23'd118;
localparam signed [DEBIT:0]  W_3_x483 = - 23'd169;
localparam signed [DEBIT:0]  W_3_x484 = - 23'd213;
localparam signed [DEBIT:0]  W_3_x485 = - 23'd246;
localparam signed [DEBIT:0]  W_3_x486 = - 23'd408;
localparam signed [DEBIT:0]  W_3_x487 = - 23'd568;
localparam signed [DEBIT:0]  W_3_x488 = - 23'd531;
localparam signed [DEBIT:0]  W_3_x489 = - 23'd378;
localparam signed [DEBIT:0]  W_3_x490 = - 23'd486;
localparam signed [DEBIT:0]  W_3_x491 = - 23'd529;
localparam signed [DEBIT:0]  W_3_x492 = - 23'd299;
localparam signed [DEBIT:0]  W_3_x493 = - 23'd84;
localparam signed [DEBIT:0]  W_3_x494 =  23'd82;
localparam signed [DEBIT:0]  W_3_x495 =  23'd20;
localparam signed [DEBIT:0]  W_3_x496 =  23'd165;
localparam signed [DEBIT:0]  W_3_x497 =  23'd112;
localparam signed [DEBIT:0]  W_3_x498 =  23'd256;
localparam signed [DEBIT:0]  W_3_x499 =  23'd226;
localparam signed [DEBIT:0]  W_3_x500 =  23'd155;
localparam signed [DEBIT:0]  W_3_x501 =  23'd264;
localparam signed [DEBIT:0]  W_3_x502 =  23'd672;
localparam signed [DEBIT:0]  W_3_x503 =  23'd914;
localparam signed [DEBIT:0]  W_3_x504 =  23'd963;
localparam signed [DEBIT:0]  W_3_x505 =  23'd960;
localparam signed [DEBIT:0]  W_3_x506 =  23'd956;
localparam signed [DEBIT:0]  W_3_x507 =  23'd976;
localparam signed [DEBIT:0]  W_3_x508 =  23'd1033;
localparam signed [DEBIT:0]  W_3_x509 =  23'd748;
localparam signed [DEBIT:0]  W_3_x510 =  23'd195;
localparam signed [DEBIT:0]  W_3_x511 =  23'd8;
localparam signed [DEBIT:0]  W_3_x512 = - 23'd3;
localparam signed [DEBIT:0]  W_3_x513 = - 23'd66;
localparam signed [DEBIT:0]  W_3_x514 = - 23'd342;
localparam signed [DEBIT:0]  W_3_x515 = - 23'd548;
localparam signed [DEBIT:0]  W_3_x516 = - 23'd544;
localparam signed [DEBIT:0]  W_3_x517 = - 23'd609;
localparam signed [DEBIT:0]  W_3_x518 = - 23'd614;
localparam signed [DEBIT:0]  W_3_x519 = - 23'd582;
localparam signed [DEBIT:0]  W_3_x520 = - 23'd275;
localparam signed [DEBIT:0]  W_3_x521 =  23'd44;
localparam signed [DEBIT:0]  W_3_x522 =  23'd44;
localparam signed [DEBIT:0]  W_3_x523 =  23'd59;
localparam signed [DEBIT:0]  W_3_x524 =  23'd180;
localparam signed [DEBIT:0]  W_3_x525 =  23'd153;
localparam signed [DEBIT:0]  W_3_x526 =  23'd202;
localparam signed [DEBIT:0]  W_3_x527 =  23'd26;
localparam signed [DEBIT:0]  W_3_x528 = - 23'd28;
localparam signed [DEBIT:0]  W_3_x529 =  23'd217;
localparam signed [DEBIT:0]  W_3_x530 =  23'd688;
localparam signed [DEBIT:0]  W_3_x531 =  23'd909;
localparam signed [DEBIT:0]  W_3_x532 =  23'd966;
localparam signed [DEBIT:0]  W_3_x533 =  23'd970;
localparam signed [DEBIT:0]  W_3_x534 =  23'd968;
localparam signed [DEBIT:0]  W_3_x535 =  23'd966;
localparam signed [DEBIT:0]  W_3_x536 =  23'd998;
localparam signed [DEBIT:0]  W_3_x537 =  23'd771;
localparam signed [DEBIT:0]  W_3_x538 =  23'd359;
localparam signed [DEBIT:0]  W_3_x539 = - 23'd5;
localparam signed [DEBIT:0]  W_3_x540 =  23'd50;
localparam signed [DEBIT:0]  W_3_x541 =  23'd8;
localparam signed [DEBIT:0]  W_3_x542 = - 23'd198;
localparam signed [DEBIT:0]  W_3_x543 = - 23'd287;
localparam signed [DEBIT:0]  W_3_x544 = - 23'd441;
localparam signed [DEBIT:0]  W_3_x545 = - 23'd448;
localparam signed [DEBIT:0]  W_3_x546 = - 23'd470;
localparam signed [DEBIT:0]  W_3_x547 = - 23'd448;
localparam signed [DEBIT:0]  W_3_x548 = - 23'd267;
localparam signed [DEBIT:0]  W_3_x549 = - 23'd61;
localparam signed [DEBIT:0]  W_3_x550 = - 23'd54;
localparam signed [DEBIT:0]  W_3_x551 = - 23'd84;
localparam signed [DEBIT:0]  W_3_x552 = - 23'd42;
localparam signed [DEBIT:0]  W_3_x553 = - 23'd2;
localparam signed [DEBIT:0]  W_3_x554 = - 23'd133;
localparam signed [DEBIT:0]  W_3_x555 = - 23'd244;
localparam signed [DEBIT:0]  W_3_x556 = - 23'd162;
localparam signed [DEBIT:0]  W_3_x557 =  23'd290;
localparam signed [DEBIT:0]  W_3_x558 =  23'd705;
localparam signed [DEBIT:0]  W_3_x559 =  23'd924;
localparam signed [DEBIT:0]  W_3_x560 =  23'd964;
localparam signed [DEBIT:0]  W_3_x561 =  23'd962;
localparam signed [DEBIT:0]  W_3_x562 =  23'd967;
localparam signed [DEBIT:0]  W_3_x563 =  23'd946;
localparam signed [DEBIT:0]  W_3_x564 =  23'd952;
localparam signed [DEBIT:0]  W_3_x565 =  23'd680;
localparam signed [DEBIT:0]  W_3_x566 =  23'd317;
localparam signed [DEBIT:0]  W_3_x567 =  23'd5;
localparam signed [DEBIT:0]  W_3_x568 = - 23'd36;
localparam signed [DEBIT:0]  W_3_x569 = - 23'd2;
localparam signed [DEBIT:0]  W_3_x570 = - 23'd27;
localparam signed [DEBIT:0]  W_3_x571 = - 23'd95;
localparam signed [DEBIT:0]  W_3_x572 = - 23'd152;
localparam signed [DEBIT:0]  W_3_x573 = - 23'd171;
localparam signed [DEBIT:0]  W_3_x574 = - 23'd228;
localparam signed [DEBIT:0]  W_3_x575 = - 23'd221;
localparam signed [DEBIT:0]  W_3_x576 = - 23'd169;
localparam signed [DEBIT:0]  W_3_x577 = - 23'd5;
localparam signed [DEBIT:0]  W_3_x578 = - 23'd46;
localparam signed [DEBIT:0]  W_3_x579 = - 23'd19;
localparam signed [DEBIT:0]  W_3_x580 = - 23'd66;
localparam signed [DEBIT:0]  W_3_x581 = - 23'd204;
localparam signed [DEBIT:0]  W_3_x582 = - 23'd288;
localparam signed [DEBIT:0]  W_3_x583 = - 23'd354;
localparam signed [DEBIT:0]  W_3_x584 = - 23'd89;
localparam signed [DEBIT:0]  W_3_x585 =  23'd366;
localparam signed [DEBIT:0]  W_3_x586 =  23'd771;
localparam signed [DEBIT:0]  W_3_x587 =  23'd934;
localparam signed [DEBIT:0]  W_3_x588 =  23'd961;
localparam signed [DEBIT:0]  W_3_x589 =  23'd973;
localparam signed [DEBIT:0]  W_3_x590 =  23'd965;
localparam signed [DEBIT:0]  W_3_x591 =  23'd941;
localparam signed [DEBIT:0]  W_3_x592 =  23'd910;
localparam signed [DEBIT:0]  W_3_x593 =  23'd631;
localparam signed [DEBIT:0]  W_3_x594 =  23'd231;
localparam signed [DEBIT:0]  W_3_x595 = - 23'd66;
localparam signed [DEBIT:0]  W_3_x596 = - 23'd165;
localparam signed [DEBIT:0]  W_3_x597 = - 23'd67;
localparam signed [DEBIT:0]  W_3_x598 = - 23'd3;
localparam signed [DEBIT:0]  W_3_x599 =  23'd38;
localparam signed [DEBIT:0]  W_3_x600 =  23'd66;
localparam signed [DEBIT:0]  W_3_x601 =  23'd29;
localparam signed [DEBIT:0]  W_3_x602 =  23'd27;
localparam signed [DEBIT:0]  W_3_x603 = - 23'd34;
localparam signed [DEBIT:0]  W_3_x604 =  23'd27;
localparam signed [DEBIT:0]  W_3_x605 =  23'd10;
localparam signed [DEBIT:0]  W_3_x606 = - 23'd52;
localparam signed [DEBIT:0]  W_3_x607 =  23'd28;
localparam signed [DEBIT:0]  W_3_x608 = - 23'd66;
localparam signed [DEBIT:0]  W_3_x609 = - 23'd289;
localparam signed [DEBIT:0]  W_3_x610 = - 23'd380;
localparam signed [DEBIT:0]  W_3_x611 = - 23'd220;
localparam signed [DEBIT:0]  W_3_x612 =  23'd183;
localparam signed [DEBIT:0]  W_3_x613 =  23'd536;
localparam signed [DEBIT:0]  W_3_x614 =  23'd866;
localparam signed [DEBIT:0]  W_3_x615 =  23'd944;
localparam signed [DEBIT:0]  W_3_x616 =  23'd957;
localparam signed [DEBIT:0]  W_3_x617 =  23'd961;
localparam signed [DEBIT:0]  W_3_x618 =  23'd963;
localparam signed [DEBIT:0]  W_3_x619 =  23'd951;
localparam signed [DEBIT:0]  W_3_x620 =  23'd937;
localparam signed [DEBIT:0]  W_3_x621 =  23'd732;
localparam signed [DEBIT:0]  W_3_x622 =  23'd308;
localparam signed [DEBIT:0]  W_3_x623 =  23'd56;
localparam signed [DEBIT:0]  W_3_x624 = - 23'd42;
localparam signed [DEBIT:0]  W_3_x625 = - 23'd119;
localparam signed [DEBIT:0]  W_3_x626 =  23'd46;
localparam signed [DEBIT:0]  W_3_x627 =  23'd132;
localparam signed [DEBIT:0]  W_3_x628 =  23'd106;
localparam signed [DEBIT:0]  W_3_x629 =  23'd88;
localparam signed [DEBIT:0]  W_3_x630 =  23'd11;
localparam signed [DEBIT:0]  W_3_x631 =  23'd10;
localparam signed [DEBIT:0]  W_3_x632 =  23'd26;
localparam signed [DEBIT:0]  W_3_x633 = - 23'd72;
localparam signed [DEBIT:0]  W_3_x634 =  23'd46;
localparam signed [DEBIT:0]  W_3_x635 =  23'd40;
localparam signed [DEBIT:0]  W_3_x636 = - 23'd105;
localparam signed [DEBIT:0]  W_3_x637 = - 23'd247;
localparam signed [DEBIT:0]  W_3_x638 = - 23'd188;
localparam signed [DEBIT:0]  W_3_x639 =  23'd107;
localparam signed [DEBIT:0]  W_3_x640 =  23'd493;
localparam signed [DEBIT:0]  W_3_x641 =  23'd744;
localparam signed [DEBIT:0]  W_3_x642 =  23'd913;
localparam signed [DEBIT:0]  W_3_x643 =  23'd965;
localparam signed [DEBIT:0]  W_3_x644 =  23'd954;
localparam signed [DEBIT:0]  W_3_x645 =  23'd965;
localparam signed [DEBIT:0]  W_3_x646 =  23'd961;
localparam signed [DEBIT:0]  W_3_x647 =  23'd969;
localparam signed [DEBIT:0]  W_3_x648 =  23'd979;
localparam signed [DEBIT:0]  W_3_x649 =  23'd927;
localparam signed [DEBIT:0]  W_3_x650 =  23'd685;
localparam signed [DEBIT:0]  W_3_x651 =  23'd406;
localparam signed [DEBIT:0]  W_3_x652 =  23'd269;
localparam signed [DEBIT:0]  W_3_x653 =  23'd106;
localparam signed [DEBIT:0]  W_3_x654 =  23'd179;
localparam signed [DEBIT:0]  W_3_x655 =  23'd130;
localparam signed [DEBIT:0]  W_3_x656 =  23'd192;
localparam signed [DEBIT:0]  W_3_x657 =  23'd222;
localparam signed [DEBIT:0]  W_3_x658 =  23'd108;
localparam signed [DEBIT:0]  W_3_x659 =  23'd48;
localparam signed [DEBIT:0]  W_3_x660 =  23'd72;
localparam signed [DEBIT:0]  W_3_x661 =  23'd100;
localparam signed [DEBIT:0]  W_3_x662 =  23'd135;
localparam signed [DEBIT:0]  W_3_x663 =  23'd55;
localparam signed [DEBIT:0]  W_3_x664 = - 23'd47;
localparam signed [DEBIT:0]  W_3_x665 = - 23'd45;
localparam signed [DEBIT:0]  W_3_x666 =  23'd179;
localparam signed [DEBIT:0]  W_3_x667 =  23'd476;
localparam signed [DEBIT:0]  W_3_x668 =  23'd737;
localparam signed [DEBIT:0]  W_3_x669 =  23'd922;
localparam signed [DEBIT:0]  W_3_x670 =  23'd955;
localparam signed [DEBIT:0]  W_3_x671 =  23'd961;
localparam signed [DEBIT:0]  W_3_x672 =  23'd963;
localparam signed [DEBIT:0]  W_3_x673 =  23'd970;
localparam signed [DEBIT:0]  W_3_x674 =  23'd959;
localparam signed [DEBIT:0]  W_3_x675 =  23'd956;
localparam signed [DEBIT:0]  W_3_x676 =  23'd1001;
localparam signed [DEBIT:0]  W_3_x677 =  23'd991;
localparam signed [DEBIT:0]  W_3_x678 =  23'd916;
localparam signed [DEBIT:0]  W_3_x679 =  23'd796;
localparam signed [DEBIT:0]  W_3_x680 =  23'd683;
localparam signed [DEBIT:0]  W_3_x681 =  23'd547;
localparam signed [DEBIT:0]  W_3_x682 =  23'd340;
localparam signed [DEBIT:0]  W_3_x683 =  23'd175;
localparam signed [DEBIT:0]  W_3_x684 =  23'd180;
localparam signed [DEBIT:0]  W_3_x685 =  23'd161;
localparam signed [DEBIT:0]  W_3_x686 =  23'd175;
localparam signed [DEBIT:0]  W_3_x687 =  23'd144;
localparam signed [DEBIT:0]  W_3_x688 =  23'd105;
localparam signed [DEBIT:0]  W_3_x689 =  23'd77;
localparam signed [DEBIT:0]  W_3_x690 =  23'd34;
localparam signed [DEBIT:0]  W_3_x691 =  23'd56;
localparam signed [DEBIT:0]  W_3_x692 =  23'd186;
localparam signed [DEBIT:0]  W_3_x693 =  23'd321;
localparam signed [DEBIT:0]  W_3_x694 =  23'd531;
localparam signed [DEBIT:0]  W_3_x695 =  23'd740;
localparam signed [DEBIT:0]  W_3_x696 =  23'd880;
localparam signed [DEBIT:0]  W_3_x697 =  23'd942;
localparam signed [DEBIT:0]  W_3_x698 =  23'd961;
localparam signed [DEBIT:0]  W_3_x699 =  23'd965;
localparam signed [DEBIT:0]  W_3_x700 =  23'd968;
localparam signed [DEBIT:0]  W_3_x701 =  23'd966;
localparam signed [DEBIT:0]  W_3_x702 =  23'd958;
localparam signed [DEBIT:0]  W_3_x703 =  23'd958;
localparam signed [DEBIT:0]  W_3_x704 =  23'd958;
localparam signed [DEBIT:0]  W_3_x705 =  23'd956;
localparam signed [DEBIT:0]  W_3_x706 =  23'd944;
localparam signed [DEBIT:0]  W_3_x707 =  23'd920;
localparam signed [DEBIT:0]  W_3_x708 =  23'd858;
localparam signed [DEBIT:0]  W_3_x709 =  23'd775;
localparam signed [DEBIT:0]  W_3_x710 =  23'd610;
localparam signed [DEBIT:0]  W_3_x711 =  23'd498;
localparam signed [DEBIT:0]  W_3_x712 =  23'd509;
localparam signed [DEBIT:0]  W_3_x713 =  23'd436;
localparam signed [DEBIT:0]  W_3_x714 =  23'd338;
localparam signed [DEBIT:0]  W_3_x715 =  23'd270;
localparam signed [DEBIT:0]  W_3_x716 =  23'd238;
localparam signed [DEBIT:0]  W_3_x717 =  23'd218;
localparam signed [DEBIT:0]  W_3_x718 =  23'd279;
localparam signed [DEBIT:0]  W_3_x719 =  23'd396;
localparam signed [DEBIT:0]  W_3_x720 =  23'd583;
localparam signed [DEBIT:0]  W_3_x721 =  23'd664;
localparam signed [DEBIT:0]  W_3_x722 =  23'd778;
localparam signed [DEBIT:0]  W_3_x723 =  23'd878;
localparam signed [DEBIT:0]  W_3_x724 =  23'd933;
localparam signed [DEBIT:0]  W_3_x725 =  23'd968;
localparam signed [DEBIT:0]  W_3_x726 =  23'd961;
localparam signed [DEBIT:0]  W_3_x727 =  23'd960;
localparam signed [DEBIT:0]  W_3_x728 =  23'd968;
localparam signed [DEBIT:0]  W_3_x729 =  23'd963;
localparam signed [DEBIT:0]  W_3_x730 =  23'd963;
localparam signed [DEBIT:0]  W_3_x731 =  23'd968;
localparam signed [DEBIT:0]  W_3_x732 =  23'd955;
localparam signed [DEBIT:0]  W_3_x733 =  23'd959;
localparam signed [DEBIT:0]  W_3_x734 =  23'd944;
localparam signed [DEBIT:0]  W_3_x735 =  23'd915;
localparam signed [DEBIT:0]  W_3_x736 =  23'd890;
localparam signed [DEBIT:0]  W_3_x737 =  23'd859;
localparam signed [DEBIT:0]  W_3_x738 =  23'd783;
localparam signed [DEBIT:0]  W_3_x739 =  23'd720;
localparam signed [DEBIT:0]  W_3_x740 =  23'd713;
localparam signed [DEBIT:0]  W_3_x741 =  23'd655;
localparam signed [DEBIT:0]  W_3_x742 =  23'd557;
localparam signed [DEBIT:0]  W_3_x743 =  23'd527;
localparam signed [DEBIT:0]  W_3_x744 =  23'd533;
localparam signed [DEBIT:0]  W_3_x745 =  23'd537;
localparam signed [DEBIT:0]  W_3_x746 =  23'd587;
localparam signed [DEBIT:0]  W_3_x747 =  23'd641;
localparam signed [DEBIT:0]  W_3_x748 =  23'd747;
localparam signed [DEBIT:0]  W_3_x749 =  23'd834;
localparam signed [DEBIT:0]  W_3_x750 =  23'd877;
localparam signed [DEBIT:0]  W_3_x751 =  23'd923;
localparam signed [DEBIT:0]  W_3_x752 =  23'd950;
localparam signed [DEBIT:0]  W_3_x753 =  23'd967;
localparam signed [DEBIT:0]  W_3_x754 =  23'd967;
localparam signed [DEBIT:0]  W_3_x755 =  23'd965;
localparam signed [DEBIT:0]  W_3_x756 =  23'd965;
localparam signed [DEBIT:0]  W_3_x757 =  23'd960;
localparam signed [DEBIT:0]  W_3_x758 =  23'd959;
localparam signed [DEBIT:0]  W_3_x759 =  23'd958;
localparam signed [DEBIT:0]  W_3_x760 =  23'd969;
localparam signed [DEBIT:0]  W_3_x761 =  23'd960;
localparam signed [DEBIT:0]  W_3_x762 =  23'd954;
localparam signed [DEBIT:0]  W_3_x763 =  23'd947;
localparam signed [DEBIT:0]  W_3_x764 =  23'd945;
localparam signed [DEBIT:0]  W_3_x765 =  23'd956;
localparam signed [DEBIT:0]  W_3_x766 =  23'd960;
localparam signed [DEBIT:0]  W_3_x767 =  23'd955;
localparam signed [DEBIT:0]  W_3_x768 =  23'd932;
localparam signed [DEBIT:0]  W_3_x769 =  23'd914;
localparam signed [DEBIT:0]  W_3_x770 =  23'd910;
localparam signed [DEBIT:0]  W_3_x771 =  23'd906;
localparam signed [DEBIT:0]  W_3_x772 =  23'd874;
localparam signed [DEBIT:0]  W_3_x773 =  23'd851;
localparam signed [DEBIT:0]  W_3_x774 =  23'd854;
localparam signed [DEBIT:0]  W_3_x775 =  23'd867;
localparam signed [DEBIT:0]  W_3_x776 =  23'd899;
localparam signed [DEBIT:0]  W_3_x777 =  23'd932;
localparam signed [DEBIT:0]  W_3_x778 =  23'd932;
localparam signed [DEBIT:0]  W_3_x779 =  23'd960;
localparam signed [DEBIT:0]  W_3_x780 =  23'd959;
localparam signed [DEBIT:0]  W_3_x781 =  23'd959;
localparam signed [DEBIT:0]  W_3_x782 =  23'd961;
localparam signed [DEBIT:0]  W_3_x783 =  23'd964;
localparam signed [DEBIT:0]  W_3_x784 =  23'd963;
localparam signed [DEBIT:0]  W_4_x1 =  23'd971;
localparam signed [DEBIT:0]  W_4_x2 =  23'd974;
localparam signed [DEBIT:0]  W_4_x3 =  23'd977;
localparam signed [DEBIT:0]  W_4_x4 =  23'd966;
localparam signed [DEBIT:0]  W_4_x5 =  23'd976;
localparam signed [DEBIT:0]  W_4_x6 =  23'd977;
localparam signed [DEBIT:0]  W_4_x7 =  23'd965;
localparam signed [DEBIT:0]  W_4_x8 =  23'd977;
localparam signed [DEBIT:0]  W_4_x9 =  23'd983;
localparam signed [DEBIT:0]  W_4_x10 =  23'd967;
localparam signed [DEBIT:0]  W_4_x11 =  23'd974;
localparam signed [DEBIT:0]  W_4_x12 =  23'd978;
localparam signed [DEBIT:0]  W_4_x13 =  23'd977;
localparam signed [DEBIT:0]  W_4_x14 =  23'd955;
localparam signed [DEBIT:0]  W_4_x15 =  23'd975;
localparam signed [DEBIT:0]  W_4_x16 =  23'd979;
localparam signed [DEBIT:0]  W_4_x17 =  23'd980;
localparam signed [DEBIT:0]  W_4_x18 =  23'd973;
localparam signed [DEBIT:0]  W_4_x19 =  23'd979;
localparam signed [DEBIT:0]  W_4_x20 =  23'd977;
localparam signed [DEBIT:0]  W_4_x21 =  23'd979;
localparam signed [DEBIT:0]  W_4_x22 =  23'd968;
localparam signed [DEBIT:0]  W_4_x23 =  23'd977;
localparam signed [DEBIT:0]  W_4_x24 =  23'd971;
localparam signed [DEBIT:0]  W_4_x25 =  23'd989;
localparam signed [DEBIT:0]  W_4_x26 =  23'd975;
localparam signed [DEBIT:0]  W_4_x27 =  23'd980;
localparam signed [DEBIT:0]  W_4_x28 =  23'd975;
localparam signed [DEBIT:0]  W_4_x29 =  23'd973;
localparam signed [DEBIT:0]  W_4_x30 =  23'd983;
localparam signed [DEBIT:0]  W_4_x31 =  23'd978;
localparam signed [DEBIT:0]  W_4_x32 =  23'd973;
localparam signed [DEBIT:0]  W_4_x33 =  23'd968;
localparam signed [DEBIT:0]  W_4_x34 =  23'd972;
localparam signed [DEBIT:0]  W_4_x35 =  23'd952;
localparam signed [DEBIT:0]  W_4_x36 =  23'd935;
localparam signed [DEBIT:0]  W_4_x37 =  23'd928;
localparam signed [DEBIT:0]  W_4_x38 =  23'd924;
localparam signed [DEBIT:0]  W_4_x39 =  23'd926;
localparam signed [DEBIT:0]  W_4_x40 =  23'd922;
localparam signed [DEBIT:0]  W_4_x41 =  23'd915;
localparam signed [DEBIT:0]  W_4_x42 =  23'd894;
localparam signed [DEBIT:0]  W_4_x43 =  23'd898;
localparam signed [DEBIT:0]  W_4_x44 =  23'd909;
localparam signed [DEBIT:0]  W_4_x45 =  23'd908;
localparam signed [DEBIT:0]  W_4_x46 =  23'd925;
localparam signed [DEBIT:0]  W_4_x47 =  23'd934;
localparam signed [DEBIT:0]  W_4_x48 =  23'd942;
localparam signed [DEBIT:0]  W_4_x49 =  23'd958;
localparam signed [DEBIT:0]  W_4_x50 =  23'd976;
localparam signed [DEBIT:0]  W_4_x51 =  23'd977;
localparam signed [DEBIT:0]  W_4_x52 =  23'd974;
localparam signed [DEBIT:0]  W_4_x53 =  23'd972;
localparam signed [DEBIT:0]  W_4_x54 =  23'd970;
localparam signed [DEBIT:0]  W_4_x55 =  23'd980;
localparam signed [DEBIT:0]  W_4_x56 =  23'd968;
localparam signed [DEBIT:0]  W_4_x57 =  23'd966;
localparam signed [DEBIT:0]  W_4_x58 =  23'd976;
localparam signed [DEBIT:0]  W_4_x59 =  23'd985;
localparam signed [DEBIT:0]  W_4_x60 =  23'd971;
localparam signed [DEBIT:0]  W_4_x61 =  23'd978;
localparam signed [DEBIT:0]  W_4_x62 =  23'd981;
localparam signed [DEBIT:0]  W_4_x63 =  23'd951;
localparam signed [DEBIT:0]  W_4_x64 =  23'd916;
localparam signed [DEBIT:0]  W_4_x65 =  23'd842;
localparam signed [DEBIT:0]  W_4_x66 =  23'd803;
localparam signed [DEBIT:0]  W_4_x67 =  23'd735;
localparam signed [DEBIT:0]  W_4_x68 =  23'd698;
localparam signed [DEBIT:0]  W_4_x69 =  23'd634;
localparam signed [DEBIT:0]  W_4_x70 =  23'd574;
localparam signed [DEBIT:0]  W_4_x71 =  23'd540;
localparam signed [DEBIT:0]  W_4_x72 =  23'd576;
localparam signed [DEBIT:0]  W_4_x73 =  23'd611;
localparam signed [DEBIT:0]  W_4_x74 =  23'd716;
localparam signed [DEBIT:0]  W_4_x75 =  23'd826;
localparam signed [DEBIT:0]  W_4_x76 =  23'd906;
localparam signed [DEBIT:0]  W_4_x77 =  23'd935;
localparam signed [DEBIT:0]  W_4_x78 =  23'd935;
localparam signed [DEBIT:0]  W_4_x79 =  23'd948;
localparam signed [DEBIT:0]  W_4_x80 =  23'd962;
localparam signed [DEBIT:0]  W_4_x81 =  23'd968;
localparam signed [DEBIT:0]  W_4_x82 =  23'd969;
localparam signed [DEBIT:0]  W_4_x83 =  23'd983;
localparam signed [DEBIT:0]  W_4_x84 =  23'd980;
localparam signed [DEBIT:0]  W_4_x85 =  23'd975;
localparam signed [DEBIT:0]  W_4_x86 =  23'd987;
localparam signed [DEBIT:0]  W_4_x87 =  23'd972;
localparam signed [DEBIT:0]  W_4_x88 =  23'd972;
localparam signed [DEBIT:0]  W_4_x89 =  23'd976;
localparam signed [DEBIT:0]  W_4_x90 =  23'd952;
localparam signed [DEBIT:0]  W_4_x91 =  23'd914;
localparam signed [DEBIT:0]  W_4_x92 =  23'd821;
localparam signed [DEBIT:0]  W_4_x93 =  23'd701;
localparam signed [DEBIT:0]  W_4_x94 =  23'd592;
localparam signed [DEBIT:0]  W_4_x95 =  23'd452;
localparam signed [DEBIT:0]  W_4_x96 =  23'd306;
localparam signed [DEBIT:0]  W_4_x97 =  23'd212;
localparam signed [DEBIT:0]  W_4_x98 =  23'd176;
localparam signed [DEBIT:0]  W_4_x99 =  23'd136;
localparam signed [DEBIT:0]  W_4_x100 =  23'd150;
localparam signed [DEBIT:0]  W_4_x101 =  23'd193;
localparam signed [DEBIT:0]  W_4_x102 =  23'd297;
localparam signed [DEBIT:0]  W_4_x103 =  23'd463;
localparam signed [DEBIT:0]  W_4_x104 =  23'd633;
localparam signed [DEBIT:0]  W_4_x105 =  23'd743;
localparam signed [DEBIT:0]  W_4_x106 =  23'd829;
localparam signed [DEBIT:0]  W_4_x107 =  23'd902;
localparam signed [DEBIT:0]  W_4_x108 =  23'd929;
localparam signed [DEBIT:0]  W_4_x109 =  23'd942;
localparam signed [DEBIT:0]  W_4_x110 =  23'd980;
localparam signed [DEBIT:0]  W_4_x111 =  23'd978;
localparam signed [DEBIT:0]  W_4_x112 =  23'd975;
localparam signed [DEBIT:0]  W_4_x113 =  23'd979;
localparam signed [DEBIT:0]  W_4_x114 =  23'd969;
localparam signed [DEBIT:0]  W_4_x115 =  23'd974;
localparam signed [DEBIT:0]  W_4_x116 =  23'd964;
localparam signed [DEBIT:0]  W_4_x117 =  23'd961;
localparam signed [DEBIT:0]  W_4_x118 =  23'd919;
localparam signed [DEBIT:0]  W_4_x119 =  23'd826;
localparam signed [DEBIT:0]  W_4_x120 =  23'd686;
localparam signed [DEBIT:0]  W_4_x121 =  23'd479;
localparam signed [DEBIT:0]  W_4_x122 =  23'd287;
localparam signed [DEBIT:0]  W_4_x123 =  23'd138;
localparam signed [DEBIT:0]  W_4_x124 =  23'd68;
localparam signed [DEBIT:0]  W_4_x125 = - 23'd37;
localparam signed [DEBIT:0]  W_4_x126 = - 23'd89;
localparam signed [DEBIT:0]  W_4_x127 = - 23'd120;
localparam signed [DEBIT:0]  W_4_x128 = - 23'd150;
localparam signed [DEBIT:0]  W_4_x129 = - 23'd139;
localparam signed [DEBIT:0]  W_4_x130 = - 23'd6;
localparam signed [DEBIT:0]  W_4_x131 =  23'd106;
localparam signed [DEBIT:0]  W_4_x132 =  23'd306;
localparam signed [DEBIT:0]  W_4_x133 =  23'd449;
localparam signed [DEBIT:0]  W_4_x134 =  23'd540;
localparam signed [DEBIT:0]  W_4_x135 =  23'd672;
localparam signed [DEBIT:0]  W_4_x136 =  23'd835;
localparam signed [DEBIT:0]  W_4_x137 =  23'd930;
localparam signed [DEBIT:0]  W_4_x138 =  23'd952;
localparam signed [DEBIT:0]  W_4_x139 =  23'd979;
localparam signed [DEBIT:0]  W_4_x140 =  23'd976;
localparam signed [DEBIT:0]  W_4_x141 =  23'd981;
localparam signed [DEBIT:0]  W_4_x142 =  23'd976;
localparam signed [DEBIT:0]  W_4_x143 =  23'd976;
localparam signed [DEBIT:0]  W_4_x144 =  23'd967;
localparam signed [DEBIT:0]  W_4_x145 =  23'd934;
localparam signed [DEBIT:0]  W_4_x146 =  23'd813;
localparam signed [DEBIT:0]  W_4_x147 =  23'd598;
localparam signed [DEBIT:0]  W_4_x148 =  23'd413;
localparam signed [DEBIT:0]  W_4_x149 =  23'd169;
localparam signed [DEBIT:0]  W_4_x150 =  23'd52;
localparam signed [DEBIT:0]  W_4_x151 = - 23'd48;
localparam signed [DEBIT:0]  W_4_x152 = - 23'd45;
localparam signed [DEBIT:0]  W_4_x153 = - 23'd56;
localparam signed [DEBIT:0]  W_4_x154 = - 23'd178;
localparam signed [DEBIT:0]  W_4_x155 = - 23'd79;
localparam signed [DEBIT:0]  W_4_x156 = - 23'd87;
localparam signed [DEBIT:0]  W_4_x157 =  23'd10;
localparam signed [DEBIT:0]  W_4_x158 = - 23'd17;
localparam signed [DEBIT:0]  W_4_x159 =  23'd61;
localparam signed [DEBIT:0]  W_4_x160 =  23'd180;
localparam signed [DEBIT:0]  W_4_x161 =  23'd203;
localparam signed [DEBIT:0]  W_4_x162 =  23'd229;
localparam signed [DEBIT:0]  W_4_x163 =  23'd440;
localparam signed [DEBIT:0]  W_4_x164 =  23'd668;
localparam signed [DEBIT:0]  W_4_x165 =  23'd779;
localparam signed [DEBIT:0]  W_4_x166 =  23'd895;
localparam signed [DEBIT:0]  W_4_x167 =  23'd964;
localparam signed [DEBIT:0]  W_4_x168 =  23'd968;
localparam signed [DEBIT:0]  W_4_x169 =  23'd974;
localparam signed [DEBIT:0]  W_4_x170 =  23'd980;
localparam signed [DEBIT:0]  W_4_x171 =  23'd964;
localparam signed [DEBIT:0]  W_4_x172 =  23'd923;
localparam signed [DEBIT:0]  W_4_x173 =  23'd840;
localparam signed [DEBIT:0]  W_4_x174 =  23'd633;
localparam signed [DEBIT:0]  W_4_x175 =  23'd364;
localparam signed [DEBIT:0]  W_4_x176 =  23'd128;
localparam signed [DEBIT:0]  W_4_x177 = - 23'd35;
localparam signed [DEBIT:0]  W_4_x178 = - 23'd145;
localparam signed [DEBIT:0]  W_4_x179 = - 23'd155;
localparam signed [DEBIT:0]  W_4_x180 = - 23'd98;
localparam signed [DEBIT:0]  W_4_x181 = - 23'd154;
localparam signed [DEBIT:0]  W_4_x182 = - 23'd179;
localparam signed [DEBIT:0]  W_4_x183 = - 23'd271;
localparam signed [DEBIT:0]  W_4_x184 = - 23'd297;
localparam signed [DEBIT:0]  W_4_x185 = - 23'd187;
localparam signed [DEBIT:0]  W_4_x186 = - 23'd28;
localparam signed [DEBIT:0]  W_4_x187 = - 23'd54;
localparam signed [DEBIT:0]  W_4_x188 =  23'd57;
localparam signed [DEBIT:0]  W_4_x189 =  23'd12;
localparam signed [DEBIT:0]  W_4_x190 =  23'd51;
localparam signed [DEBIT:0]  W_4_x191 =  23'd271;
localparam signed [DEBIT:0]  W_4_x192 =  23'd549;
localparam signed [DEBIT:0]  W_4_x193 =  23'd609;
localparam signed [DEBIT:0]  W_4_x194 =  23'd728;
localparam signed [DEBIT:0]  W_4_x195 =  23'd895;
localparam signed [DEBIT:0]  W_4_x196 =  23'd972;
localparam signed [DEBIT:0]  W_4_x197 =  23'd979;
localparam signed [DEBIT:0]  W_4_x198 =  23'd972;
localparam signed [DEBIT:0]  W_4_x199 =  23'd928;
localparam signed [DEBIT:0]  W_4_x200 =  23'd834;
localparam signed [DEBIT:0]  W_4_x201 =  23'd653;
localparam signed [DEBIT:0]  W_4_x202 =  23'd378;
localparam signed [DEBIT:0]  W_4_x203 =  23'd76;
localparam signed [DEBIT:0]  W_4_x204 = - 23'd104;
localparam signed [DEBIT:0]  W_4_x205 = - 23'd52;
localparam signed [DEBIT:0]  W_4_x206 = - 23'd1;
localparam signed [DEBIT:0]  W_4_x207 = - 23'd45;
localparam signed [DEBIT:0]  W_4_x208 = - 23'd206;
localparam signed [DEBIT:0]  W_4_x209 = - 23'd370;
localparam signed [DEBIT:0]  W_4_x210 = - 23'd418;
localparam signed [DEBIT:0]  W_4_x211 = - 23'd537;
localparam signed [DEBIT:0]  W_4_x212 = - 23'd690;
localparam signed [DEBIT:0]  W_4_x213 = - 23'd584;
localparam signed [DEBIT:0]  W_4_x214 = - 23'd285;
localparam signed [DEBIT:0]  W_4_x215 = - 23'd92;
localparam signed [DEBIT:0]  W_4_x216 = - 23'd1;
localparam signed [DEBIT:0]  W_4_x217 = - 23'd127;
localparam signed [DEBIT:0]  W_4_x218 = - 23'd86;
localparam signed [DEBIT:0]  W_4_x219 =  23'd31;
localparam signed [DEBIT:0]  W_4_x220 =  23'd286;
localparam signed [DEBIT:0]  W_4_x221 =  23'd453;
localparam signed [DEBIT:0]  W_4_x222 =  23'd671;
localparam signed [DEBIT:0]  W_4_x223 =  23'd862;
localparam signed [DEBIT:0]  W_4_x224 =  23'd961;
localparam signed [DEBIT:0]  W_4_x225 =  23'd966;
localparam signed [DEBIT:0]  W_4_x226 =  23'd911;
localparam signed [DEBIT:0]  W_4_x227 =  23'd842;
localparam signed [DEBIT:0]  W_4_x228 =  23'd650;
localparam signed [DEBIT:0]  W_4_x229 =  23'd407;
localparam signed [DEBIT:0]  W_4_x230 =  23'd129;
localparam signed [DEBIT:0]  W_4_x231 = - 23'd134;
localparam signed [DEBIT:0]  W_4_x232 = - 23'd184;
localparam signed [DEBIT:0]  W_4_x233 = - 23'd97;
localparam signed [DEBIT:0]  W_4_x234 =  23'd69;
localparam signed [DEBIT:0]  W_4_x235 = - 23'd146;
localparam signed [DEBIT:0]  W_4_x236 = - 23'd290;
localparam signed [DEBIT:0]  W_4_x237 = - 23'd483;
localparam signed [DEBIT:0]  W_4_x238 = - 23'd512;
localparam signed [DEBIT:0]  W_4_x239 = - 23'd671;
localparam signed [DEBIT:0]  W_4_x240 = - 23'd747;
localparam signed [DEBIT:0]  W_4_x241 = - 23'd495;
localparam signed [DEBIT:0]  W_4_x242 = - 23'd356;
localparam signed [DEBIT:0]  W_4_x243 = - 23'd251;
localparam signed [DEBIT:0]  W_4_x244 = - 23'd65;
localparam signed [DEBIT:0]  W_4_x245 = - 23'd138;
localparam signed [DEBIT:0]  W_4_x246 = - 23'd238;
localparam signed [DEBIT:0]  W_4_x247 = - 23'd57;
localparam signed [DEBIT:0]  W_4_x248 =  23'd224;
localparam signed [DEBIT:0]  W_4_x249 =  23'd431;
localparam signed [DEBIT:0]  W_4_x250 =  23'd664;
localparam signed [DEBIT:0]  W_4_x251 =  23'd869;
localparam signed [DEBIT:0]  W_4_x252 =  23'd956;
localparam signed [DEBIT:0]  W_4_x253 =  23'd969;
localparam signed [DEBIT:0]  W_4_x254 =  23'd911;
localparam signed [DEBIT:0]  W_4_x255 =  23'd809;
localparam signed [DEBIT:0]  W_4_x256 =  23'd588;
localparam signed [DEBIT:0]  W_4_x257 =  23'd320;
localparam signed [DEBIT:0]  W_4_x258 = - 23'd23;
localparam signed [DEBIT:0]  W_4_x259 = - 23'd353;
localparam signed [DEBIT:0]  W_4_x260 = - 23'd258;
localparam signed [DEBIT:0]  W_4_x261 = - 23'd174;
localparam signed [DEBIT:0]  W_4_x262 = - 23'd137;
localparam signed [DEBIT:0]  W_4_x263 = - 23'd286;
localparam signed [DEBIT:0]  W_4_x264 = - 23'd348;
localparam signed [DEBIT:0]  W_4_x265 = - 23'd268;
localparam signed [DEBIT:0]  W_4_x266 = - 23'd436;
localparam signed [DEBIT:0]  W_4_x267 = - 23'd849;
localparam signed [DEBIT:0]  W_4_x268 = - 23'd552;
localparam signed [DEBIT:0]  W_4_x269 = - 23'd199;
localparam signed [DEBIT:0]  W_4_x270 = - 23'd186;
localparam signed [DEBIT:0]  W_4_x271 = - 23'd159;
localparam signed [DEBIT:0]  W_4_x272 = - 23'd95;
localparam signed [DEBIT:0]  W_4_x273 = - 23'd165;
localparam signed [DEBIT:0]  W_4_x274 = - 23'd254;
localparam signed [DEBIT:0]  W_4_x275 = - 23'd129;
localparam signed [DEBIT:0]  W_4_x276 =  23'd154;
localparam signed [DEBIT:0]  W_4_x277 =  23'd445;
localparam signed [DEBIT:0]  W_4_x278 =  23'd692;
localparam signed [DEBIT:0]  W_4_x279 =  23'd872;
localparam signed [DEBIT:0]  W_4_x280 =  23'd962;
localparam signed [DEBIT:0]  W_4_x281 =  23'd973;
localparam signed [DEBIT:0]  W_4_x282 =  23'd918;
localparam signed [DEBIT:0]  W_4_x283 =  23'd810;
localparam signed [DEBIT:0]  W_4_x284 =  23'd596;
localparam signed [DEBIT:0]  W_4_x285 =  23'd283;
localparam signed [DEBIT:0]  W_4_x286 = - 23'd124;
localparam signed [DEBIT:0]  W_4_x287 = - 23'd423;
localparam signed [DEBIT:0]  W_4_x288 = - 23'd303;
localparam signed [DEBIT:0]  W_4_x289 = - 23'd158;
localparam signed [DEBIT:0]  W_4_x290 = - 23'd102;
localparam signed [DEBIT:0]  W_4_x291 = - 23'd207;
localparam signed [DEBIT:0]  W_4_x292 = - 23'd139;
localparam signed [DEBIT:0]  W_4_x293 =  23'd26;
localparam signed [DEBIT:0]  W_4_x294 = - 23'd409;
localparam signed [DEBIT:0]  W_4_x295 = - 23'd868;
localparam signed [DEBIT:0]  W_4_x296 = - 23'd366;
localparam signed [DEBIT:0]  W_4_x297 = - 23'd93;
localparam signed [DEBIT:0]  W_4_x298 = - 23'd71;
localparam signed [DEBIT:0]  W_4_x299 = - 23'd126;
localparam signed [DEBIT:0]  W_4_x300 = - 23'd54;
localparam signed [DEBIT:0]  W_4_x301 = - 23'd214;
localparam signed [DEBIT:0]  W_4_x302 = - 23'd347;
localparam signed [DEBIT:0]  W_4_x303 = - 23'd188;
localparam signed [DEBIT:0]  W_4_x304 =  23'd116;
localparam signed [DEBIT:0]  W_4_x305 =  23'd523;
localparam signed [DEBIT:0]  W_4_x306 =  23'd753;
localparam signed [DEBIT:0]  W_4_x307 =  23'd907;
localparam signed [DEBIT:0]  W_4_x308 =  23'd967;
localparam signed [DEBIT:0]  W_4_x309 =  23'd968;
localparam signed [DEBIT:0]  W_4_x310 =  23'd938;
localparam signed [DEBIT:0]  W_4_x311 =  23'd819;
localparam signed [DEBIT:0]  W_4_x312 =  23'd604;
localparam signed [DEBIT:0]  W_4_x313 =  23'd285;
localparam signed [DEBIT:0]  W_4_x314 = - 23'd143;
localparam signed [DEBIT:0]  W_4_x315 = - 23'd374;
localparam signed [DEBIT:0]  W_4_x316 = - 23'd290;
localparam signed [DEBIT:0]  W_4_x317 = - 23'd14;
localparam signed [DEBIT:0]  W_4_x318 = - 23'd24;
localparam signed [DEBIT:0]  W_4_x319 =  23'd78;
localparam signed [DEBIT:0]  W_4_x320 =  23'd312;
localparam signed [DEBIT:0]  W_4_x321 =  23'd263;
localparam signed [DEBIT:0]  W_4_x322 = - 23'd442;
localparam signed [DEBIT:0]  W_4_x323 = - 23'd664;
localparam signed [DEBIT:0]  W_4_x324 = - 23'd24;
localparam signed [DEBIT:0]  W_4_x325 =  23'd257;
localparam signed [DEBIT:0]  W_4_x326 =  23'd63;
localparam signed [DEBIT:0]  W_4_x327 = - 23'd98;
localparam signed [DEBIT:0]  W_4_x328 = - 23'd95;
localparam signed [DEBIT:0]  W_4_x329 = - 23'd286;
localparam signed [DEBIT:0]  W_4_x330 = - 23'd313;
localparam signed [DEBIT:0]  W_4_x331 = - 23'd177;
localparam signed [DEBIT:0]  W_4_x332 =  23'd153;
localparam signed [DEBIT:0]  W_4_x333 =  23'd585;
localparam signed [DEBIT:0]  W_4_x334 =  23'd848;
localparam signed [DEBIT:0]  W_4_x335 =  23'd938;
localparam signed [DEBIT:0]  W_4_x336 =  23'd967;
localparam signed [DEBIT:0]  W_4_x337 =  23'd971;
localparam signed [DEBIT:0]  W_4_x338 =  23'd939;
localparam signed [DEBIT:0]  W_4_x339 =  23'd861;
localparam signed [DEBIT:0]  W_4_x340 =  23'd687;
localparam signed [DEBIT:0]  W_4_x341 =  23'd355;
localparam signed [DEBIT:0]  W_4_x342 = - 23'd44;
localparam signed [DEBIT:0]  W_4_x343 = - 23'd256;
localparam signed [DEBIT:0]  W_4_x344 = - 23'd20;
localparam signed [DEBIT:0]  W_4_x345 =  23'd220;
localparam signed [DEBIT:0]  W_4_x346 =  23'd179;
localparam signed [DEBIT:0]  W_4_x347 =  23'd282;
localparam signed [DEBIT:0]  W_4_x348 =  23'd588;
localparam signed [DEBIT:0]  W_4_x349 =  23'd378;
localparam signed [DEBIT:0]  W_4_x350 = - 23'd259;
localparam signed [DEBIT:0]  W_4_x351 = - 23'd413;
localparam signed [DEBIT:0]  W_4_x352 =  23'd86;
localparam signed [DEBIT:0]  W_4_x353 =  23'd298;
localparam signed [DEBIT:0]  W_4_x354 =  23'd83;
localparam signed [DEBIT:0]  W_4_x355 = - 23'd12;
localparam signed [DEBIT:0]  W_4_x356 = - 23'd52;
localparam signed [DEBIT:0]  W_4_x357 = - 23'd322;
localparam signed [DEBIT:0]  W_4_x358 = - 23'd294;
localparam signed [DEBIT:0]  W_4_x359 = - 23'd136;
localparam signed [DEBIT:0]  W_4_x360 =  23'd181;
localparam signed [DEBIT:0]  W_4_x361 =  23'd556;
localparam signed [DEBIT:0]  W_4_x362 =  23'd879;
localparam signed [DEBIT:0]  W_4_x363 =  23'd958;
localparam signed [DEBIT:0]  W_4_x364 =  23'd971;
localparam signed [DEBIT:0]  W_4_x365 =  23'd970;
localparam signed [DEBIT:0]  W_4_x366 =  23'd963;
localparam signed [DEBIT:0]  W_4_x367 =  23'd928;
localparam signed [DEBIT:0]  W_4_x368 =  23'd780;
localparam signed [DEBIT:0]  W_4_x369 =  23'd501;
localparam signed [DEBIT:0]  W_4_x370 =  23'd155;
localparam signed [DEBIT:0]  W_4_x371 =  23'd55;
localparam signed [DEBIT:0]  W_4_x372 =  23'd317;
localparam signed [DEBIT:0]  W_4_x373 =  23'd355;
localparam signed [DEBIT:0]  W_4_x374 =  23'd275;
localparam signed [DEBIT:0]  W_4_x375 =  23'd438;
localparam signed [DEBIT:0]  W_4_x376 =  23'd589;
localparam signed [DEBIT:0]  W_4_x377 =  23'd304;
localparam signed [DEBIT:0]  W_4_x378 = - 23'd174;
localparam signed [DEBIT:0]  W_4_x379 = - 23'd194;
localparam signed [DEBIT:0]  W_4_x380 =  23'd95;
localparam signed [DEBIT:0]  W_4_x381 =  23'd162;
localparam signed [DEBIT:0]  W_4_x382 =  23'd157;
localparam signed [DEBIT:0]  W_4_x383 =  23'd3;
localparam signed [DEBIT:0]  W_4_x384 =  23'd56;
localparam signed [DEBIT:0]  W_4_x385 = - 23'd68;
localparam signed [DEBIT:0]  W_4_x386 = - 23'd92;
localparam signed [DEBIT:0]  W_4_x387 = - 23'd32;
localparam signed [DEBIT:0]  W_4_x388 =  23'd163;
localparam signed [DEBIT:0]  W_4_x389 =  23'd502;
localparam signed [DEBIT:0]  W_4_x390 =  23'd874;
localparam signed [DEBIT:0]  W_4_x391 =  23'd961;
localparam signed [DEBIT:0]  W_4_x392 =  23'd956;
localparam signed [DEBIT:0]  W_4_x393 =  23'd987;
localparam signed [DEBIT:0]  W_4_x394 =  23'd973;
localparam signed [DEBIT:0]  W_4_x395 =  23'd957;
localparam signed [DEBIT:0]  W_4_x396 =  23'd862;
localparam signed [DEBIT:0]  W_4_x397 =  23'd661;
localparam signed [DEBIT:0]  W_4_x398 =  23'd331;
localparam signed [DEBIT:0]  W_4_x399 =  23'd261;
localparam signed [DEBIT:0]  W_4_x400 =  23'd410;
localparam signed [DEBIT:0]  W_4_x401 =  23'd250;
localparam signed [DEBIT:0]  W_4_x402 =  23'd167;
localparam signed [DEBIT:0]  W_4_x403 =  23'd247;
localparam signed [DEBIT:0]  W_4_x404 =  23'd419;
localparam signed [DEBIT:0]  W_4_x405 =  23'd204;
localparam signed [DEBIT:0]  W_4_x406 = - 23'd97;
localparam signed [DEBIT:0]  W_4_x407 = - 23'd76;
localparam signed [DEBIT:0]  W_4_x408 =  23'd29;
localparam signed [DEBIT:0]  W_4_x409 =  23'd134;
localparam signed [DEBIT:0]  W_4_x410 =  23'd181;
localparam signed [DEBIT:0]  W_4_x411 =  23'd98;
localparam signed [DEBIT:0]  W_4_x412 =  23'd277;
localparam signed [DEBIT:0]  W_4_x413 =  23'd182;
localparam signed [DEBIT:0]  W_4_x414 =  23'd11;
localparam signed [DEBIT:0]  W_4_x415 = - 23'd3;
localparam signed [DEBIT:0]  W_4_x416 =  23'd123;
localparam signed [DEBIT:0]  W_4_x417 =  23'd434;
localparam signed [DEBIT:0]  W_4_x418 =  23'd828;
localparam signed [DEBIT:0]  W_4_x419 =  23'd946;
localparam signed [DEBIT:0]  W_4_x420 =  23'd972;
localparam signed [DEBIT:0]  W_4_x421 =  23'd972;
localparam signed [DEBIT:0]  W_4_x422 =  23'd971;
localparam signed [DEBIT:0]  W_4_x423 =  23'd973;
localparam signed [DEBIT:0]  W_4_x424 =  23'd872;
localparam signed [DEBIT:0]  W_4_x425 =  23'd669;
localparam signed [DEBIT:0]  W_4_x426 =  23'd300;
localparam signed [DEBIT:0]  W_4_x427 =  23'd232;
localparam signed [DEBIT:0]  W_4_x428 =  23'd299;
localparam signed [DEBIT:0]  W_4_x429 =  23'd219;
localparam signed [DEBIT:0]  W_4_x430 =  23'd141;
localparam signed [DEBIT:0]  W_4_x431 =  23'd40;
localparam signed [DEBIT:0]  W_4_x432 =  23'd210;
localparam signed [DEBIT:0]  W_4_x433 =  23'd180;
localparam signed [DEBIT:0]  W_4_x434 = - 23'd4;
localparam signed [DEBIT:0]  W_4_x435 =  23'd54;
localparam signed [DEBIT:0]  W_4_x436 =  23'd259;
localparam signed [DEBIT:0]  W_4_x437 =  23'd290;
localparam signed [DEBIT:0]  W_4_x438 =  23'd193;
localparam signed [DEBIT:0]  W_4_x439 =  23'd180;
localparam signed [DEBIT:0]  W_4_x440 =  23'd295;
localparam signed [DEBIT:0]  W_4_x441 =  23'd129;
localparam signed [DEBIT:0]  W_4_x442 = - 23'd22;
localparam signed [DEBIT:0]  W_4_x443 = - 23'd29;
localparam signed [DEBIT:0]  W_4_x444 =  23'd63;
localparam signed [DEBIT:0]  W_4_x445 =  23'd347;
localparam signed [DEBIT:0]  W_4_x446 =  23'd729;
localparam signed [DEBIT:0]  W_4_x447 =  23'd935;
localparam signed [DEBIT:0]  W_4_x448 =  23'd970;
localparam signed [DEBIT:0]  W_4_x449 =  23'd970;
localparam signed [DEBIT:0]  W_4_x450 =  23'd979;
localparam signed [DEBIT:0]  W_4_x451 =  23'd974;
localparam signed [DEBIT:0]  W_4_x452 =  23'd807;
localparam signed [DEBIT:0]  W_4_x453 =  23'd521;
localparam signed [DEBIT:0]  W_4_x454 =  23'd222;
localparam signed [DEBIT:0]  W_4_x455 =  23'd154;
localparam signed [DEBIT:0]  W_4_x456 =  23'd306;
localparam signed [DEBIT:0]  W_4_x457 =  23'd356;
localparam signed [DEBIT:0]  W_4_x458 =  23'd132;
localparam signed [DEBIT:0]  W_4_x459 =  23'd27;
localparam signed [DEBIT:0]  W_4_x460 =  23'd22;
localparam signed [DEBIT:0]  W_4_x461 =  23'd104;
localparam signed [DEBIT:0]  W_4_x462 =  23'd75;
localparam signed [DEBIT:0]  W_4_x463 =  23'd302;
localparam signed [DEBIT:0]  W_4_x464 =  23'd394;
localparam signed [DEBIT:0]  W_4_x465 =  23'd283;
localparam signed [DEBIT:0]  W_4_x466 =  23'd329;
localparam signed [DEBIT:0]  W_4_x467 =  23'd312;
localparam signed [DEBIT:0]  W_4_x468 =  23'd197;
localparam signed [DEBIT:0]  W_4_x469 =  23'd89;
localparam signed [DEBIT:0]  W_4_x470 = - 23'd117;
localparam signed [DEBIT:0]  W_4_x471 = - 23'd108;
localparam signed [DEBIT:0]  W_4_x472 = - 23'd3;
localparam signed [DEBIT:0]  W_4_x473 =  23'd272;
localparam signed [DEBIT:0]  W_4_x474 =  23'd680;
localparam signed [DEBIT:0]  W_4_x475 =  23'd915;
localparam signed [DEBIT:0]  W_4_x476 =  23'd966;
localparam signed [DEBIT:0]  W_4_x477 =  23'd977;
localparam signed [DEBIT:0]  W_4_x478 =  23'd980;
localparam signed [DEBIT:0]  W_4_x479 =  23'd960;
localparam signed [DEBIT:0]  W_4_x480 =  23'd746;
localparam signed [DEBIT:0]  W_4_x481 =  23'd411;
localparam signed [DEBIT:0]  W_4_x482 =  23'd83;
localparam signed [DEBIT:0]  W_4_x483 =  23'd114;
localparam signed [DEBIT:0]  W_4_x484 =  23'd275;
localparam signed [DEBIT:0]  W_4_x485 =  23'd354;
localparam signed [DEBIT:0]  W_4_x486 =  23'd264;
localparam signed [DEBIT:0]  W_4_x487 =  23'd29;
localparam signed [DEBIT:0]  W_4_x488 = - 23'd49;
localparam signed [DEBIT:0]  W_4_x489 =  23'd198;
localparam signed [DEBIT:0]  W_4_x490 =  23'd373;
localparam signed [DEBIT:0]  W_4_x491 =  23'd546;
localparam signed [DEBIT:0]  W_4_x492 =  23'd383;
localparam signed [DEBIT:0]  W_4_x493 =  23'd192;
localparam signed [DEBIT:0]  W_4_x494 =  23'd156;
localparam signed [DEBIT:0]  W_4_x495 =  23'd110;
localparam signed [DEBIT:0]  W_4_x496 = - 23'd62;
localparam signed [DEBIT:0]  W_4_x497 = - 23'd248;
localparam signed [DEBIT:0]  W_4_x498 = - 23'd401;
localparam signed [DEBIT:0]  W_4_x499 = - 23'd333;
localparam signed [DEBIT:0]  W_4_x500 = - 23'd46;
localparam signed [DEBIT:0]  W_4_x501 =  23'd296;
localparam signed [DEBIT:0]  W_4_x502 =  23'd732;
localparam signed [DEBIT:0]  W_4_x503 =  23'd939;
localparam signed [DEBIT:0]  W_4_x504 =  23'd969;
localparam signed [DEBIT:0]  W_4_x505 =  23'd970;
localparam signed [DEBIT:0]  W_4_x506 =  23'd982;
localparam signed [DEBIT:0]  W_4_x507 =  23'd960;
localparam signed [DEBIT:0]  W_4_x508 =  23'd690;
localparam signed [DEBIT:0]  W_4_x509 =  23'd324;
localparam signed [DEBIT:0]  W_4_x510 = - 23'd15;
localparam signed [DEBIT:0]  W_4_x511 = - 23'd17;
localparam signed [DEBIT:0]  W_4_x512 =  23'd86;
localparam signed [DEBIT:0]  W_4_x513 =  23'd147;
localparam signed [DEBIT:0]  W_4_x514 =  23'd80;
localparam signed [DEBIT:0]  W_4_x515 = - 23'd226;
localparam signed [DEBIT:0]  W_4_x516 = - 23'd218;
localparam signed [DEBIT:0]  W_4_x517 =  23'd0;
localparam signed [DEBIT:0]  W_4_x518 =  23'd167;
localparam signed [DEBIT:0]  W_4_x519 =  23'd227;
localparam signed [DEBIT:0]  W_4_x520 =  23'd51;
localparam signed [DEBIT:0]  W_4_x521 = - 23'd54;
localparam signed [DEBIT:0]  W_4_x522 = - 23'd311;
localparam signed [DEBIT:0]  W_4_x523 = - 23'd354;
localparam signed [DEBIT:0]  W_4_x524 = - 23'd361;
localparam signed [DEBIT:0]  W_4_x525 = - 23'd449;
localparam signed [DEBIT:0]  W_4_x526 = - 23'd585;
localparam signed [DEBIT:0]  W_4_x527 = - 23'd512;
localparam signed [DEBIT:0]  W_4_x528 = - 23'd71;
localparam signed [DEBIT:0]  W_4_x529 =  23'd448;
localparam signed [DEBIT:0]  W_4_x530 =  23'd795;
localparam signed [DEBIT:0]  W_4_x531 =  23'd955;
localparam signed [DEBIT:0]  W_4_x532 =  23'd976;
localparam signed [DEBIT:0]  W_4_x533 =  23'd977;
localparam signed [DEBIT:0]  W_4_x534 =  23'd970;
localparam signed [DEBIT:0]  W_4_x535 =  23'd947;
localparam signed [DEBIT:0]  W_4_x536 =  23'd656;
localparam signed [DEBIT:0]  W_4_x537 =  23'd261;
localparam signed [DEBIT:0]  W_4_x538 = - 23'd41;
localparam signed [DEBIT:0]  W_4_x539 = - 23'd270;
localparam signed [DEBIT:0]  W_4_x540 = - 23'd324;
localparam signed [DEBIT:0]  W_4_x541 = - 23'd408;
localparam signed [DEBIT:0]  W_4_x542 = - 23'd510;
localparam signed [DEBIT:0]  W_4_x543 = - 23'd648;
localparam signed [DEBIT:0]  W_4_x544 = - 23'd638;
localparam signed [DEBIT:0]  W_4_x545 = - 23'd493;
localparam signed [DEBIT:0]  W_4_x546 = - 23'd319;
localparam signed [DEBIT:0]  W_4_x547 = - 23'd201;
localparam signed [DEBIT:0]  W_4_x548 = - 23'd246;
localparam signed [DEBIT:0]  W_4_x549 = - 23'd282;
localparam signed [DEBIT:0]  W_4_x550 = - 23'd537;
localparam signed [DEBIT:0]  W_4_x551 = - 23'd536;
localparam signed [DEBIT:0]  W_4_x552 = - 23'd587;
localparam signed [DEBIT:0]  W_4_x553 = - 23'd584;
localparam signed [DEBIT:0]  W_4_x554 = - 23'd662;
localparam signed [DEBIT:0]  W_4_x555 = - 23'd533;
localparam signed [DEBIT:0]  W_4_x556 =  23'd37;
localparam signed [DEBIT:0]  W_4_x557 =  23'd620;
localparam signed [DEBIT:0]  W_4_x558 =  23'd869;
localparam signed [DEBIT:0]  W_4_x559 =  23'd949;
localparam signed [DEBIT:0]  W_4_x560 =  23'd982;
localparam signed [DEBIT:0]  W_4_x561 =  23'd967;
localparam signed [DEBIT:0]  W_4_x562 =  23'd971;
localparam signed [DEBIT:0]  W_4_x563 =  23'd925;
localparam signed [DEBIT:0]  W_4_x564 =  23'd665;
localparam signed [DEBIT:0]  W_4_x565 =  23'd221;
localparam signed [DEBIT:0]  W_4_x566 = - 23'd28;
localparam signed [DEBIT:0]  W_4_x567 = - 23'd336;
localparam signed [DEBIT:0]  W_4_x568 = - 23'd514;
localparam signed [DEBIT:0]  W_4_x569 = - 23'd647;
localparam signed [DEBIT:0]  W_4_x570 = - 23'd648;
localparam signed [DEBIT:0]  W_4_x571 = - 23'd567;
localparam signed [DEBIT:0]  W_4_x572 = - 23'd528;
localparam signed [DEBIT:0]  W_4_x573 = - 23'd455;
localparam signed [DEBIT:0]  W_4_x574 = - 23'd513;
localparam signed [DEBIT:0]  W_4_x575 = - 23'd415;
localparam signed [DEBIT:0]  W_4_x576 = - 23'd348;
localparam signed [DEBIT:0]  W_4_x577 = - 23'd247;
localparam signed [DEBIT:0]  W_4_x578 = - 23'd337;
localparam signed [DEBIT:0]  W_4_x579 = - 23'd367;
localparam signed [DEBIT:0]  W_4_x580 = - 23'd500;
localparam signed [DEBIT:0]  W_4_x581 = - 23'd581;
localparam signed [DEBIT:0]  W_4_x582 = - 23'd521;
localparam signed [DEBIT:0]  W_4_x583 = - 23'd314;
localparam signed [DEBIT:0]  W_4_x584 =  23'd230;
localparam signed [DEBIT:0]  W_4_x585 =  23'd714;
localparam signed [DEBIT:0]  W_4_x586 =  23'd904;
localparam signed [DEBIT:0]  W_4_x587 =  23'd961;
localparam signed [DEBIT:0]  W_4_x588 =  23'd972;
localparam signed [DEBIT:0]  W_4_x589 =  23'd972;
localparam signed [DEBIT:0]  W_4_x590 =  23'd969;
localparam signed [DEBIT:0]  W_4_x591 =  23'd932;
localparam signed [DEBIT:0]  W_4_x592 =  23'd742;
localparam signed [DEBIT:0]  W_4_x593 =  23'd361;
localparam signed [DEBIT:0]  W_4_x594 = - 23'd1;
localparam signed [DEBIT:0]  W_4_x595 = - 23'd344;
localparam signed [DEBIT:0]  W_4_x596 = - 23'd604;
localparam signed [DEBIT:0]  W_4_x597 = - 23'd569;
localparam signed [DEBIT:0]  W_4_x598 = - 23'd476;
localparam signed [DEBIT:0]  W_4_x599 = - 23'd258;
localparam signed [DEBIT:0]  W_4_x600 = - 23'd54;
localparam signed [DEBIT:0]  W_4_x601 = - 23'd124;
localparam signed [DEBIT:0]  W_4_x602 = - 23'd115;
localparam signed [DEBIT:0]  W_4_x603 = - 23'd123;
localparam signed [DEBIT:0]  W_4_x604 =  23'd8;
localparam signed [DEBIT:0]  W_4_x605 = - 23'd95;
localparam signed [DEBIT:0]  W_4_x606 = - 23'd43;
localparam signed [DEBIT:0]  W_4_x607 = - 23'd49;
localparam signed [DEBIT:0]  W_4_x608 = - 23'd147;
localparam signed [DEBIT:0]  W_4_x609 = - 23'd292;
localparam signed [DEBIT:0]  W_4_x610 = - 23'd237;
localparam signed [DEBIT:0]  W_4_x611 =  23'd3;
localparam signed [DEBIT:0]  W_4_x612 =  23'd459;
localparam signed [DEBIT:0]  W_4_x613 =  23'd775;
localparam signed [DEBIT:0]  W_4_x614 =  23'd925;
localparam signed [DEBIT:0]  W_4_x615 =  23'd962;
localparam signed [DEBIT:0]  W_4_x616 =  23'd968;
localparam signed [DEBIT:0]  W_4_x617 =  23'd972;
localparam signed [DEBIT:0]  W_4_x618 =  23'd973;
localparam signed [DEBIT:0]  W_4_x619 =  23'd941;
localparam signed [DEBIT:0]  W_4_x620 =  23'd830;
localparam signed [DEBIT:0]  W_4_x621 =  23'd575;
localparam signed [DEBIT:0]  W_4_x622 =  23'd231;
localparam signed [DEBIT:0]  W_4_x623 = - 23'd119;
localparam signed [DEBIT:0]  W_4_x624 = - 23'd392;
localparam signed [DEBIT:0]  W_4_x625 = - 23'd401;
localparam signed [DEBIT:0]  W_4_x626 = - 23'd278;
localparam signed [DEBIT:0]  W_4_x627 = - 23'd70;
localparam signed [DEBIT:0]  W_4_x628 =  23'd4;
localparam signed [DEBIT:0]  W_4_x629 = - 23'd15;
localparam signed [DEBIT:0]  W_4_x630 =  23'd8;
localparam signed [DEBIT:0]  W_4_x631 = - 23'd8;
localparam signed [DEBIT:0]  W_4_x632 =  23'd164;
localparam signed [DEBIT:0]  W_4_x633 =  23'd165;
localparam signed [DEBIT:0]  W_4_x634 =  23'd237;
localparam signed [DEBIT:0]  W_4_x635 =  23'd186;
localparam signed [DEBIT:0]  W_4_x636 =  23'd104;
localparam signed [DEBIT:0]  W_4_x637 =  23'd37;
localparam signed [DEBIT:0]  W_4_x638 =  23'd87;
localparam signed [DEBIT:0]  W_4_x639 =  23'd331;
localparam signed [DEBIT:0]  W_4_x640 =  23'd689;
localparam signed [DEBIT:0]  W_4_x641 =  23'd888;
localparam signed [DEBIT:0]  W_4_x642 =  23'd948;
localparam signed [DEBIT:0]  W_4_x643 =  23'd974;
localparam signed [DEBIT:0]  W_4_x644 =  23'd978;
localparam signed [DEBIT:0]  W_4_x645 =  23'd972;
localparam signed [DEBIT:0]  W_4_x646 =  23'd977;
localparam signed [DEBIT:0]  W_4_x647 =  23'd957;
localparam signed [DEBIT:0]  W_4_x648 =  23'd909;
localparam signed [DEBIT:0]  W_4_x649 =  23'd787;
localparam signed [DEBIT:0]  W_4_x650 =  23'd565;
localparam signed [DEBIT:0]  W_4_x651 =  23'd254;
localparam signed [DEBIT:0]  W_4_x652 =  23'd25;
localparam signed [DEBIT:0]  W_4_x653 = - 23'd126;
localparam signed [DEBIT:0]  W_4_x654 = - 23'd175;
localparam signed [DEBIT:0]  W_4_x655 = - 23'd162;
localparam signed [DEBIT:0]  W_4_x656 = - 23'd103;
localparam signed [DEBIT:0]  W_4_x657 = - 23'd100;
localparam signed [DEBIT:0]  W_4_x658 = - 23'd103;
localparam signed [DEBIT:0]  W_4_x659 = - 23'd17;
localparam signed [DEBIT:0]  W_4_x660 =  23'd138;
localparam signed [DEBIT:0]  W_4_x661 =  23'd259;
localparam signed [DEBIT:0]  W_4_x662 =  23'd351;
localparam signed [DEBIT:0]  W_4_x663 =  23'd309;
localparam signed [DEBIT:0]  W_4_x664 =  23'd360;
localparam signed [DEBIT:0]  W_4_x665 =  23'd371;
localparam signed [DEBIT:0]  W_4_x666 =  23'd438;
localparam signed [DEBIT:0]  W_4_x667 =  23'd636;
localparam signed [DEBIT:0]  W_4_x668 =  23'd852;
localparam signed [DEBIT:0]  W_4_x669 =  23'd954;
localparam signed [DEBIT:0]  W_4_x670 =  23'd971;
localparam signed [DEBIT:0]  W_4_x671 =  23'd983;
localparam signed [DEBIT:0]  W_4_x672 =  23'd973;
localparam signed [DEBIT:0]  W_4_x673 =  23'd975;
localparam signed [DEBIT:0]  W_4_x674 =  23'd984;
localparam signed [DEBIT:0]  W_4_x675 =  23'd980;
localparam signed [DEBIT:0]  W_4_x676 =  23'd963;
localparam signed [DEBIT:0]  W_4_x677 =  23'd918;
localparam signed [DEBIT:0]  W_4_x678 =  23'd811;
localparam signed [DEBIT:0]  W_4_x679 =  23'd691;
localparam signed [DEBIT:0]  W_4_x680 =  23'd458;
localparam signed [DEBIT:0]  W_4_x681 =  23'd275;
localparam signed [DEBIT:0]  W_4_x682 =  23'd137;
localparam signed [DEBIT:0]  W_4_x683 =  23'd53;
localparam signed [DEBIT:0]  W_4_x684 =  23'd96;
localparam signed [DEBIT:0]  W_4_x685 =  23'd66;
localparam signed [DEBIT:0]  W_4_x686 =  23'd32;
localparam signed [DEBIT:0]  W_4_x687 =  23'd66;
localparam signed [DEBIT:0]  W_4_x688 =  23'd54;
localparam signed [DEBIT:0]  W_4_x689 =  23'd135;
localparam signed [DEBIT:0]  W_4_x690 =  23'd113;
localparam signed [DEBIT:0]  W_4_x691 =  23'd250;
localparam signed [DEBIT:0]  W_4_x692 =  23'd410;
localparam signed [DEBIT:0]  W_4_x693 =  23'd485;
localparam signed [DEBIT:0]  W_4_x694 =  23'd579;
localparam signed [DEBIT:0]  W_4_x695 =  23'd750;
localparam signed [DEBIT:0]  W_4_x696 =  23'd887;
localparam signed [DEBIT:0]  W_4_x697 =  23'd963;
localparam signed [DEBIT:0]  W_4_x698 =  23'd970;
localparam signed [DEBIT:0]  W_4_x699 =  23'd986;
localparam signed [DEBIT:0]  W_4_x700 =  23'd984;
localparam signed [DEBIT:0]  W_4_x701 =  23'd975;
localparam signed [DEBIT:0]  W_4_x702 =  23'd967;
localparam signed [DEBIT:0]  W_4_x703 =  23'd960;
localparam signed [DEBIT:0]  W_4_x704 =  23'd979;
localparam signed [DEBIT:0]  W_4_x705 =  23'd956;
localparam signed [DEBIT:0]  W_4_x706 =  23'd952;
localparam signed [DEBIT:0]  W_4_x707 =  23'd884;
localparam signed [DEBIT:0]  W_4_x708 =  23'd771;
localparam signed [DEBIT:0]  W_4_x709 =  23'd622;
localparam signed [DEBIT:0]  W_4_x710 =  23'd495;
localparam signed [DEBIT:0]  W_4_x711 =  23'd348;
localparam signed [DEBIT:0]  W_4_x712 =  23'd224;
localparam signed [DEBIT:0]  W_4_x713 =  23'd130;
localparam signed [DEBIT:0]  W_4_x714 =  23'd132;
localparam signed [DEBIT:0]  W_4_x715 =  23'd142;
localparam signed [DEBIT:0]  W_4_x716 =  23'd136;
localparam signed [DEBIT:0]  W_4_x717 =  23'd60;
localparam signed [DEBIT:0]  W_4_x718 =  23'd83;
localparam signed [DEBIT:0]  W_4_x719 =  23'd236;
localparam signed [DEBIT:0]  W_4_x720 =  23'd394;
localparam signed [DEBIT:0]  W_4_x721 =  23'd560;
localparam signed [DEBIT:0]  W_4_x722 =  23'd706;
localparam signed [DEBIT:0]  W_4_x723 =  23'd818;
localparam signed [DEBIT:0]  W_4_x724 =  23'd934;
localparam signed [DEBIT:0]  W_4_x725 =  23'd967;
localparam signed [DEBIT:0]  W_4_x726 =  23'd974;
localparam signed [DEBIT:0]  W_4_x727 =  23'd974;
localparam signed [DEBIT:0]  W_4_x728 =  23'd974;
localparam signed [DEBIT:0]  W_4_x729 =  23'd981;
localparam signed [DEBIT:0]  W_4_x730 =  23'd976;
localparam signed [DEBIT:0]  W_4_x731 =  23'd980;
localparam signed [DEBIT:0]  W_4_x732 =  23'd980;
localparam signed [DEBIT:0]  W_4_x733 =  23'd979;
localparam signed [DEBIT:0]  W_4_x734 =  23'd971;
localparam signed [DEBIT:0]  W_4_x735 =  23'd895;
localparam signed [DEBIT:0]  W_4_x736 =  23'd848;
localparam signed [DEBIT:0]  W_4_x737 =  23'd787;
localparam signed [DEBIT:0]  W_4_x738 =  23'd723;
localparam signed [DEBIT:0]  W_4_x739 =  23'd647;
localparam signed [DEBIT:0]  W_4_x740 =  23'd579;
localparam signed [DEBIT:0]  W_4_x741 =  23'd566;
localparam signed [DEBIT:0]  W_4_x742 =  23'd514;
localparam signed [DEBIT:0]  W_4_x743 =  23'd466;
localparam signed [DEBIT:0]  W_4_x744 =  23'd456;
localparam signed [DEBIT:0]  W_4_x745 =  23'd415;
localparam signed [DEBIT:0]  W_4_x746 =  23'd443;
localparam signed [DEBIT:0]  W_4_x747 =  23'd536;
localparam signed [DEBIT:0]  W_4_x748 =  23'd627;
localparam signed [DEBIT:0]  W_4_x749 =  23'd766;
localparam signed [DEBIT:0]  W_4_x750 =  23'd861;
localparam signed [DEBIT:0]  W_4_x751 =  23'd914;
localparam signed [DEBIT:0]  W_4_x752 =  23'd958;
localparam signed [DEBIT:0]  W_4_x753 =  23'd975;
localparam signed [DEBIT:0]  W_4_x754 =  23'd980;
localparam signed [DEBIT:0]  W_4_x755 =  23'd986;
localparam signed [DEBIT:0]  W_4_x756 =  23'd974;
localparam signed [DEBIT:0]  W_4_x757 =  23'd973;
localparam signed [DEBIT:0]  W_4_x758 =  23'd972;
localparam signed [DEBIT:0]  W_4_x759 =  23'd975;
localparam signed [DEBIT:0]  W_4_x760 =  23'd967;
localparam signed [DEBIT:0]  W_4_x761 =  23'd976;
localparam signed [DEBIT:0]  W_4_x762 =  23'd978;
localparam signed [DEBIT:0]  W_4_x763 =  23'd954;
localparam signed [DEBIT:0]  W_4_x764 =  23'd942;
localparam signed [DEBIT:0]  W_4_x765 =  23'd944;
localparam signed [DEBIT:0]  W_4_x766 =  23'd959;
localparam signed [DEBIT:0]  W_4_x767 =  23'd961;
localparam signed [DEBIT:0]  W_4_x768 =  23'd926;
localparam signed [DEBIT:0]  W_4_x769 =  23'd896;
localparam signed [DEBIT:0]  W_4_x770 =  23'd889;
localparam signed [DEBIT:0]  W_4_x771 =  23'd850;
localparam signed [DEBIT:0]  W_4_x772 =  23'd877;
localparam signed [DEBIT:0]  W_4_x773 =  23'd860;
localparam signed [DEBIT:0]  W_4_x774 =  23'd867;
localparam signed [DEBIT:0]  W_4_x775 =  23'd863;
localparam signed [DEBIT:0]  W_4_x776 =  23'd902;
localparam signed [DEBIT:0]  W_4_x777 =  23'd944;
localparam signed [DEBIT:0]  W_4_x778 =  23'd950;
localparam signed [DEBIT:0]  W_4_x779 =  23'd960;
localparam signed [DEBIT:0]  W_4_x780 =  23'd977;
localparam signed [DEBIT:0]  W_4_x781 =  23'd972;
localparam signed [DEBIT:0]  W_4_x782 =  23'd972;
localparam signed [DEBIT:0]  W_4_x783 =  23'd979;
localparam signed [DEBIT:0]  W_4_x784 =  23'd971;
localparam signed [DEBIT:0]  W_5_x1 =  23'd975;
localparam signed [DEBIT:0]  W_5_x2 =  23'd983;
localparam signed [DEBIT:0]  W_5_x3 =  23'd979;
localparam signed [DEBIT:0]  W_5_x4 =  23'd977;
localparam signed [DEBIT:0]  W_5_x5 =  23'd979;
localparam signed [DEBIT:0]  W_5_x6 =  23'd983;
localparam signed [DEBIT:0]  W_5_x7 =  23'd971;
localparam signed [DEBIT:0]  W_5_x8 =  23'd975;
localparam signed [DEBIT:0]  W_5_x9 =  23'd975;
localparam signed [DEBIT:0]  W_5_x10 =  23'd968;
localparam signed [DEBIT:0]  W_5_x11 =  23'd982;
localparam signed [DEBIT:0]  W_5_x12 =  23'd974;
localparam signed [DEBIT:0]  W_5_x13 =  23'd977;
localparam signed [DEBIT:0]  W_5_x14 =  23'd970;
localparam signed [DEBIT:0]  W_5_x15 =  23'd982;
localparam signed [DEBIT:0]  W_5_x16 =  23'd984;
localparam signed [DEBIT:0]  W_5_x17 =  23'd981;
localparam signed [DEBIT:0]  W_5_x18 =  23'd977;
localparam signed [DEBIT:0]  W_5_x19 =  23'd979;
localparam signed [DEBIT:0]  W_5_x20 =  23'd975;
localparam signed [DEBIT:0]  W_5_x21 =  23'd973;
localparam signed [DEBIT:0]  W_5_x22 =  23'd976;
localparam signed [DEBIT:0]  W_5_x23 =  23'd980;
localparam signed [DEBIT:0]  W_5_x24 =  23'd977;
localparam signed [DEBIT:0]  W_5_x25 =  23'd975;
localparam signed [DEBIT:0]  W_5_x26 =  23'd972;
localparam signed [DEBIT:0]  W_5_x27 =  23'd969;
localparam signed [DEBIT:0]  W_5_x28 =  23'd982;
localparam signed [DEBIT:0]  W_5_x29 =  23'd979;
localparam signed [DEBIT:0]  W_5_x30 =  23'd978;
localparam signed [DEBIT:0]  W_5_x31 =  23'd978;
localparam signed [DEBIT:0]  W_5_x32 =  23'd978;
localparam signed [DEBIT:0]  W_5_x33 =  23'd977;
localparam signed [DEBIT:0]  W_5_x34 =  23'd986;
localparam signed [DEBIT:0]  W_5_x35 =  23'd977;
localparam signed [DEBIT:0]  W_5_x36 =  23'd973;
localparam signed [DEBIT:0]  W_5_x37 =  23'd976;
localparam signed [DEBIT:0]  W_5_x38 =  23'd964;
localparam signed [DEBIT:0]  W_5_x39 =  23'd955;
localparam signed [DEBIT:0]  W_5_x40 =  23'd970;
localparam signed [DEBIT:0]  W_5_x41 =  23'd963;
localparam signed [DEBIT:0]  W_5_x42 =  23'd964;
localparam signed [DEBIT:0]  W_5_x43 =  23'd958;
localparam signed [DEBIT:0]  W_5_x44 =  23'd964;
localparam signed [DEBIT:0]  W_5_x45 =  23'd964;
localparam signed [DEBIT:0]  W_5_x46 =  23'd981;
localparam signed [DEBIT:0]  W_5_x47 =  23'd981;
localparam signed [DEBIT:0]  W_5_x48 =  23'd977;
localparam signed [DEBIT:0]  W_5_x49 =  23'd976;
localparam signed [DEBIT:0]  W_5_x50 =  23'd970;
localparam signed [DEBIT:0]  W_5_x51 =  23'd975;
localparam signed [DEBIT:0]  W_5_x52 =  23'd973;
localparam signed [DEBIT:0]  W_5_x53 =  23'd985;
localparam signed [DEBIT:0]  W_5_x54 =  23'd988;
localparam signed [DEBIT:0]  W_5_x55 =  23'd977;
localparam signed [DEBIT:0]  W_5_x56 =  23'd973;
localparam signed [DEBIT:0]  W_5_x57 =  23'd989;
localparam signed [DEBIT:0]  W_5_x58 =  23'd974;
localparam signed [DEBIT:0]  W_5_x59 =  23'd983;
localparam signed [DEBIT:0]  W_5_x60 =  23'd984;
localparam signed [DEBIT:0]  W_5_x61 =  23'd977;
localparam signed [DEBIT:0]  W_5_x62 =  23'd980;
localparam signed [DEBIT:0]  W_5_x63 =  23'd977;
localparam signed [DEBIT:0]  W_5_x64 =  23'd963;
localparam signed [DEBIT:0]  W_5_x65 =  23'd927;
localparam signed [DEBIT:0]  W_5_x66 =  23'd887;
localparam signed [DEBIT:0]  W_5_x67 =  23'd863;
localparam signed [DEBIT:0]  W_5_x68 =  23'd834;
localparam signed [DEBIT:0]  W_5_x69 =  23'd779;
localparam signed [DEBIT:0]  W_5_x70 =  23'd768;
localparam signed [DEBIT:0]  W_5_x71 =  23'd750;
localparam signed [DEBIT:0]  W_5_x72 =  23'd715;
localparam signed [DEBIT:0]  W_5_x73 =  23'd714;
localparam signed [DEBIT:0]  W_5_x74 =  23'd771;
localparam signed [DEBIT:0]  W_5_x75 =  23'd801;
localparam signed [DEBIT:0]  W_5_x76 =  23'd825;
localparam signed [DEBIT:0]  W_5_x77 =  23'd872;
localparam signed [DEBIT:0]  W_5_x78 =  23'd893;
localparam signed [DEBIT:0]  W_5_x79 =  23'd909;
localparam signed [DEBIT:0]  W_5_x80 =  23'd945;
localparam signed [DEBIT:0]  W_5_x81 =  23'd971;
localparam signed [DEBIT:0]  W_5_x82 =  23'd981;
localparam signed [DEBIT:0]  W_5_x83 =  23'd984;
localparam signed [DEBIT:0]  W_5_x84 =  23'd981;
localparam signed [DEBIT:0]  W_5_x85 =  23'd989;
localparam signed [DEBIT:0]  W_5_x86 =  23'd973;
localparam signed [DEBIT:0]  W_5_x87 =  23'd978;
localparam signed [DEBIT:0]  W_5_x88 =  23'd981;
localparam signed [DEBIT:0]  W_5_x89 =  23'd976;
localparam signed [DEBIT:0]  W_5_x90 =  23'd957;
localparam signed [DEBIT:0]  W_5_x91 =  23'd925;
localparam signed [DEBIT:0]  W_5_x92 =  23'd836;
localparam signed [DEBIT:0]  W_5_x93 =  23'd725;
localparam signed [DEBIT:0]  W_5_x94 =  23'd623;
localparam signed [DEBIT:0]  W_5_x95 =  23'd529;
localparam signed [DEBIT:0]  W_5_x96 =  23'd396;
localparam signed [DEBIT:0]  W_5_x97 =  23'd352;
localparam signed [DEBIT:0]  W_5_x98 =  23'd346;
localparam signed [DEBIT:0]  W_5_x99 =  23'd271;
localparam signed [DEBIT:0]  W_5_x100 =  23'd197;
localparam signed [DEBIT:0]  W_5_x101 =  23'd223;
localparam signed [DEBIT:0]  W_5_x102 =  23'd281;
localparam signed [DEBIT:0]  W_5_x103 =  23'd357;
localparam signed [DEBIT:0]  W_5_x104 =  23'd423;
localparam signed [DEBIT:0]  W_5_x105 =  23'd536;
localparam signed [DEBIT:0]  W_5_x106 =  23'd644;
localparam signed [DEBIT:0]  W_5_x107 =  23'd760;
localparam signed [DEBIT:0]  W_5_x108 =  23'd852;
localparam signed [DEBIT:0]  W_5_x109 =  23'd917;
localparam signed [DEBIT:0]  W_5_x110 =  23'd970;
localparam signed [DEBIT:0]  W_5_x111 =  23'd979;
localparam signed [DEBIT:0]  W_5_x112 =  23'd980;
localparam signed [DEBIT:0]  W_5_x113 =  23'd977;
localparam signed [DEBIT:0]  W_5_x114 =  23'd983;
localparam signed [DEBIT:0]  W_5_x115 =  23'd979;
localparam signed [DEBIT:0]  W_5_x116 =  23'd977;
localparam signed [DEBIT:0]  W_5_x117 =  23'd954;
localparam signed [DEBIT:0]  W_5_x118 =  23'd874;
localparam signed [DEBIT:0]  W_5_x119 =  23'd736;
localparam signed [DEBIT:0]  W_5_x120 =  23'd511;
localparam signed [DEBIT:0]  W_5_x121 =  23'd249;
localparam signed [DEBIT:0]  W_5_x122 =  23'd62;
localparam signed [DEBIT:0]  W_5_x123 =  23'd19;
localparam signed [DEBIT:0]  W_5_x124 = - 23'd18;
localparam signed [DEBIT:0]  W_5_x125 = - 23'd129;
localparam signed [DEBIT:0]  W_5_x126 = - 23'd133;
localparam signed [DEBIT:0]  W_5_x127 = - 23'd31;
localparam signed [DEBIT:0]  W_5_x128 =  23'd8;
localparam signed [DEBIT:0]  W_5_x129 =  23'd11;
localparam signed [DEBIT:0]  W_5_x130 =  23'd6;
localparam signed [DEBIT:0]  W_5_x131 =  23'd64;
localparam signed [DEBIT:0]  W_5_x132 =  23'd67;
localparam signed [DEBIT:0]  W_5_x133 =  23'd181;
localparam signed [DEBIT:0]  W_5_x134 =  23'd442;
localparam signed [DEBIT:0]  W_5_x135 =  23'd646;
localparam signed [DEBIT:0]  W_5_x136 =  23'd842;
localparam signed [DEBIT:0]  W_5_x137 =  23'd925;
localparam signed [DEBIT:0]  W_5_x138 =  23'd954;
localparam signed [DEBIT:0]  W_5_x139 =  23'd976;
localparam signed [DEBIT:0]  W_5_x140 =  23'd980;
localparam signed [DEBIT:0]  W_5_x141 =  23'd980;
localparam signed [DEBIT:0]  W_5_x142 =  23'd979;
localparam signed [DEBIT:0]  W_5_x143 =  23'd964;
localparam signed [DEBIT:0]  W_5_x144 =  23'd966;
localparam signed [DEBIT:0]  W_5_x145 =  23'd855;
localparam signed [DEBIT:0]  W_5_x146 =  23'd603;
localparam signed [DEBIT:0]  W_5_x147 =  23'd258;
localparam signed [DEBIT:0]  W_5_x148 = - 23'd42;
localparam signed [DEBIT:0]  W_5_x149 = - 23'd217;
localparam signed [DEBIT:0]  W_5_x150 = - 23'd241;
localparam signed [DEBIT:0]  W_5_x151 = - 23'd146;
localparam signed [DEBIT:0]  W_5_x152 = - 23'd49;
localparam signed [DEBIT:0]  W_5_x153 = - 23'd88;
localparam signed [DEBIT:0]  W_5_x154 = - 23'd245;
localparam signed [DEBIT:0]  W_5_x155 = - 23'd109;
localparam signed [DEBIT:0]  W_5_x156 = - 23'd106;
localparam signed [DEBIT:0]  W_5_x157 = - 23'd118;
localparam signed [DEBIT:0]  W_5_x158 =  23'd2;
localparam signed [DEBIT:0]  W_5_x159 = - 23'd13;
localparam signed [DEBIT:0]  W_5_x160 = - 23'd7;
localparam signed [DEBIT:0]  W_5_x161 =  23'd124;
localparam signed [DEBIT:0]  W_5_x162 =  23'd209;
localparam signed [DEBIT:0]  W_5_x163 =  23'd497;
localparam signed [DEBIT:0]  W_5_x164 =  23'd765;
localparam signed [DEBIT:0]  W_5_x165 =  23'd891;
localparam signed [DEBIT:0]  W_5_x166 =  23'd916;
localparam signed [DEBIT:0]  W_5_x167 =  23'd961;
localparam signed [DEBIT:0]  W_5_x168 =  23'd979;
localparam signed [DEBIT:0]  W_5_x169 =  23'd988;
localparam signed [DEBIT:0]  W_5_x170 =  23'd974;
localparam signed [DEBIT:0]  W_5_x171 =  23'd968;
localparam signed [DEBIT:0]  W_5_x172 =  23'd864;
localparam signed [DEBIT:0]  W_5_x173 =  23'd632;
localparam signed [DEBIT:0]  W_5_x174 =  23'd294;
localparam signed [DEBIT:0]  W_5_x175 = - 23'd54;
localparam signed [DEBIT:0]  W_5_x176 = - 23'd227;
localparam signed [DEBIT:0]  W_5_x177 = - 23'd271;
localparam signed [DEBIT:0]  W_5_x178 = - 23'd141;
localparam signed [DEBIT:0]  W_5_x179 = - 23'd57;
localparam signed [DEBIT:0]  W_5_x180 =  23'd59;
localparam signed [DEBIT:0]  W_5_x181 = - 23'd9;
localparam signed [DEBIT:0]  W_5_x182 = - 23'd89;
localparam signed [DEBIT:0]  W_5_x183 =  23'd29;
localparam signed [DEBIT:0]  W_5_x184 = - 23'd49;
localparam signed [DEBIT:0]  W_5_x185 =  23'd6;
localparam signed [DEBIT:0]  W_5_x186 =  23'd42;
localparam signed [DEBIT:0]  W_5_x187 =  23'd18;
localparam signed [DEBIT:0]  W_5_x188 =  23'd10;
localparam signed [DEBIT:0]  W_5_x189 =  23'd34;
localparam signed [DEBIT:0]  W_5_x190 = - 23'd49;
localparam signed [DEBIT:0]  W_5_x191 =  23'd213;
localparam signed [DEBIT:0]  W_5_x192 =  23'd645;
localparam signed [DEBIT:0]  W_5_x193 =  23'd909;
localparam signed [DEBIT:0]  W_5_x194 =  23'd900;
localparam signed [DEBIT:0]  W_5_x195 =  23'd936;
localparam signed [DEBIT:0]  W_5_x196 =  23'd969;
localparam signed [DEBIT:0]  W_5_x197 =  23'd981;
localparam signed [DEBIT:0]  W_5_x198 =  23'd977;
localparam signed [DEBIT:0]  W_5_x199 =  23'd931;
localparam signed [DEBIT:0]  W_5_x200 =  23'd739;
localparam signed [DEBIT:0]  W_5_x201 =  23'd395;
localparam signed [DEBIT:0]  W_5_x202 =  23'd72;
localparam signed [DEBIT:0]  W_5_x203 = - 23'd157;
localparam signed [DEBIT:0]  W_5_x204 = - 23'd123;
localparam signed [DEBIT:0]  W_5_x205 =  23'd90;
localparam signed [DEBIT:0]  W_5_x206 =  23'd101;
localparam signed [DEBIT:0]  W_5_x207 =  23'd258;
localparam signed [DEBIT:0]  W_5_x208 =  23'd248;
localparam signed [DEBIT:0]  W_5_x209 =  23'd71;
localparam signed [DEBIT:0]  W_5_x210 = - 23'd106;
localparam signed [DEBIT:0]  W_5_x211 = - 23'd108;
localparam signed [DEBIT:0]  W_5_x212 = - 23'd170;
localparam signed [DEBIT:0]  W_5_x213 = - 23'd111;
localparam signed [DEBIT:0]  W_5_x214 =  23'd63;
localparam signed [DEBIT:0]  W_5_x215 =  23'd90;
localparam signed [DEBIT:0]  W_5_x216 =  23'd66;
localparam signed [DEBIT:0]  W_5_x217 =  23'd4;
localparam signed [DEBIT:0]  W_5_x218 = - 23'd76;
localparam signed [DEBIT:0]  W_5_x219 =  23'd77;
localparam signed [DEBIT:0]  W_5_x220 =  23'd585;
localparam signed [DEBIT:0]  W_5_x221 =  23'd1031;
localparam signed [DEBIT:0]  W_5_x222 =  23'd1074;
localparam signed [DEBIT:0]  W_5_x223 =  23'd958;
localparam signed [DEBIT:0]  W_5_x224 =  23'd993;
localparam signed [DEBIT:0]  W_5_x225 =  23'd989;
localparam signed [DEBIT:0]  W_5_x226 =  23'd928;
localparam signed [DEBIT:0]  W_5_x227 =  23'd819;
localparam signed [DEBIT:0]  W_5_x228 =  23'd573;
localparam signed [DEBIT:0]  W_5_x229 =  23'd146;
localparam signed [DEBIT:0]  W_5_x230 = - 23'd75;
localparam signed [DEBIT:0]  W_5_x231 = - 23'd202;
localparam signed [DEBIT:0]  W_5_x232 = - 23'd34;
localparam signed [DEBIT:0]  W_5_x233 =  23'd139;
localparam signed [DEBIT:0]  W_5_x234 =  23'd175;
localparam signed [DEBIT:0]  W_5_x235 =  23'd136;
localparam signed [DEBIT:0]  W_5_x236 =  23'd143;
localparam signed [DEBIT:0]  W_5_x237 = - 23'd41;
localparam signed [DEBIT:0]  W_5_x238 = - 23'd232;
localparam signed [DEBIT:0]  W_5_x239 = - 23'd294;
localparam signed [DEBIT:0]  W_5_x240 = - 23'd348;
localparam signed [DEBIT:0]  W_5_x241 = - 23'd278;
localparam signed [DEBIT:0]  W_5_x242 = - 23'd118;
localparam signed [DEBIT:0]  W_5_x243 = - 23'd14;
localparam signed [DEBIT:0]  W_5_x244 =  23'd26;
localparam signed [DEBIT:0]  W_5_x245 =  23'd114;
localparam signed [DEBIT:0]  W_5_x246 =  23'd35;
localparam signed [DEBIT:0]  W_5_x247 =  23'd67;
localparam signed [DEBIT:0]  W_5_x248 =  23'd608;
localparam signed [DEBIT:0]  W_5_x249 =  23'd1264;
localparam signed [DEBIT:0]  W_5_x250 =  23'd1249;
localparam signed [DEBIT:0]  W_5_x251 =  23'd984;
localparam signed [DEBIT:0]  W_5_x252 =  23'd968;
localparam signed [DEBIT:0]  W_5_x253 =  23'd973;
localparam signed [DEBIT:0]  W_5_x254 =  23'd895;
localparam signed [DEBIT:0]  W_5_x255 =  23'd788;
localparam signed [DEBIT:0]  W_5_x256 =  23'd504;
localparam signed [DEBIT:0]  W_5_x257 =  23'd129;
localparam signed [DEBIT:0]  W_5_x258 = - 23'd78;
localparam signed [DEBIT:0]  W_5_x259 = - 23'd232;
localparam signed [DEBIT:0]  W_5_x260 = - 23'd23;
localparam signed [DEBIT:0]  W_5_x261 =  23'd111;
localparam signed [DEBIT:0]  W_5_x262 =  23'd45;
localparam signed [DEBIT:0]  W_5_x263 = - 23'd8;
localparam signed [DEBIT:0]  W_5_x264 =  23'd207;
localparam signed [DEBIT:0]  W_5_x265 =  23'd27;
localparam signed [DEBIT:0]  W_5_x266 = - 23'd194;
localparam signed [DEBIT:0]  W_5_x267 = - 23'd344;
localparam signed [DEBIT:0]  W_5_x268 = - 23'd438;
localparam signed [DEBIT:0]  W_5_x269 = - 23'd418;
localparam signed [DEBIT:0]  W_5_x270 = - 23'd271;
localparam signed [DEBIT:0]  W_5_x271 = - 23'd239;
localparam signed [DEBIT:0]  W_5_x272 = - 23'd180;
localparam signed [DEBIT:0]  W_5_x273 = - 23'd16;
localparam signed [DEBIT:0]  W_5_x274 =  23'd31;
localparam signed [DEBIT:0]  W_5_x275 =  23'd5;
localparam signed [DEBIT:0]  W_5_x276 =  23'd438;
localparam signed [DEBIT:0]  W_5_x277 =  23'd1245;
localparam signed [DEBIT:0]  W_5_x278 =  23'd1335;
localparam signed [DEBIT:0]  W_5_x279 =  23'd1025;
localparam signed [DEBIT:0]  W_5_x280 =  23'd986;
localparam signed [DEBIT:0]  W_5_x281 =  23'd986;
localparam signed [DEBIT:0]  W_5_x282 =  23'd903;
localparam signed [DEBIT:0]  W_5_x283 =  23'd760;
localparam signed [DEBIT:0]  W_5_x284 =  23'd514;
localparam signed [DEBIT:0]  W_5_x285 =  23'd205;
localparam signed [DEBIT:0]  W_5_x286 = - 23'd79;
localparam signed [DEBIT:0]  W_5_x287 = - 23'd213;
localparam signed [DEBIT:0]  W_5_x288 =  23'd12;
localparam signed [DEBIT:0]  W_5_x289 =  23'd158;
localparam signed [DEBIT:0]  W_5_x290 =  23'd144;
localparam signed [DEBIT:0]  W_5_x291 =  23'd155;
localparam signed [DEBIT:0]  W_5_x292 =  23'd318;
localparam signed [DEBIT:0]  W_5_x293 =  23'd296;
localparam signed [DEBIT:0]  W_5_x294 =  23'd200;
localparam signed [DEBIT:0]  W_5_x295 = - 23'd47;
localparam signed [DEBIT:0]  W_5_x296 = - 23'd262;
localparam signed [DEBIT:0]  W_5_x297 = - 23'd439;
localparam signed [DEBIT:0]  W_5_x298 = - 23'd473;
localparam signed [DEBIT:0]  W_5_x299 = - 23'd522;
localparam signed [DEBIT:0]  W_5_x300 = - 23'd522;
localparam signed [DEBIT:0]  W_5_x301 = - 23'd411;
localparam signed [DEBIT:0]  W_5_x302 = - 23'd311;
localparam signed [DEBIT:0]  W_5_x303 = - 23'd403;
localparam signed [DEBIT:0]  W_5_x304 = - 23'd14;
localparam signed [DEBIT:0]  W_5_x305 =  23'd826;
localparam signed [DEBIT:0]  W_5_x306 =  23'd1326;
localparam signed [DEBIT:0]  W_5_x307 =  23'd1043;
localparam signed [DEBIT:0]  W_5_x308 =  23'd975;
localparam signed [DEBIT:0]  W_5_x309 =  23'd973;
localparam signed [DEBIT:0]  W_5_x310 =  23'd915;
localparam signed [DEBIT:0]  W_5_x311 =  23'd794;
localparam signed [DEBIT:0]  W_5_x312 =  23'd564;
localparam signed [DEBIT:0]  W_5_x313 =  23'd316;
localparam signed [DEBIT:0]  W_5_x314 = - 23'd23;
localparam signed [DEBIT:0]  W_5_x315 = - 23'd168;
localparam signed [DEBIT:0]  W_5_x316 =  23'd7;
localparam signed [DEBIT:0]  W_5_x317 =  23'd220;
localparam signed [DEBIT:0]  W_5_x318 =  23'd201;
localparam signed [DEBIT:0]  W_5_x319 =  23'd225;
localparam signed [DEBIT:0]  W_5_x320 =  23'd355;
localparam signed [DEBIT:0]  W_5_x321 =  23'd348;
localparam signed [DEBIT:0]  W_5_x322 =  23'd255;
localparam signed [DEBIT:0]  W_5_x323 = - 23'd14;
localparam signed [DEBIT:0]  W_5_x324 = - 23'd77;
localparam signed [DEBIT:0]  W_5_x325 = - 23'd264;
localparam signed [DEBIT:0]  W_5_x326 = - 23'd412;
localparam signed [DEBIT:0]  W_5_x327 = - 23'd543;
localparam signed [DEBIT:0]  W_5_x328 = - 23'd757;
localparam signed [DEBIT:0]  W_5_x329 = - 23'd826;
localparam signed [DEBIT:0]  W_5_x330 = - 23'd783;
localparam signed [DEBIT:0]  W_5_x331 = - 23'd856;
localparam signed [DEBIT:0]  W_5_x332 = - 23'd511;
localparam signed [DEBIT:0]  W_5_x333 =  23'd323;
localparam signed [DEBIT:0]  W_5_x334 =  23'd1079;
localparam signed [DEBIT:0]  W_5_x335 =  23'd1003;
localparam signed [DEBIT:0]  W_5_x336 =  23'd982;
localparam signed [DEBIT:0]  W_5_x337 =  23'd986;
localparam signed [DEBIT:0]  W_5_x338 =  23'd942;
localparam signed [DEBIT:0]  W_5_x339 =  23'd841;
localparam signed [DEBIT:0]  W_5_x340 =  23'd681;
localparam signed [DEBIT:0]  W_5_x341 =  23'd435;
localparam signed [DEBIT:0]  W_5_x342 =  23'd112;
localparam signed [DEBIT:0]  W_5_x343 = - 23'd28;
localparam signed [DEBIT:0]  W_5_x344 =  23'd83;
localparam signed [DEBIT:0]  W_5_x345 =  23'd199;
localparam signed [DEBIT:0]  W_5_x346 =  23'd169;
localparam signed [DEBIT:0]  W_5_x347 =  23'd216;
localparam signed [DEBIT:0]  W_5_x348 =  23'd252;
localparam signed [DEBIT:0]  W_5_x349 =  23'd368;
localparam signed [DEBIT:0]  W_5_x350 =  23'd258;
localparam signed [DEBIT:0]  W_5_x351 = - 23'd56;
localparam signed [DEBIT:0]  W_5_x352 = - 23'd131;
localparam signed [DEBIT:0]  W_5_x353 = - 23'd247;
localparam signed [DEBIT:0]  W_5_x354 = - 23'd223;
localparam signed [DEBIT:0]  W_5_x355 = - 23'd294;
localparam signed [DEBIT:0]  W_5_x356 = - 23'd408;
localparam signed [DEBIT:0]  W_5_x357 = - 23'd582;
localparam signed [DEBIT:0]  W_5_x358 = - 23'd639;
localparam signed [DEBIT:0]  W_5_x359 = - 23'd873;
localparam signed [DEBIT:0]  W_5_x360 = - 23'd674;
localparam signed [DEBIT:0]  W_5_x361 =  23'd38;
localparam signed [DEBIT:0]  W_5_x362 =  23'd901;
localparam signed [DEBIT:0]  W_5_x363 =  23'd976;
localparam signed [DEBIT:0]  W_5_x364 =  23'd979;
localparam signed [DEBIT:0]  W_5_x365 =  23'd976;
localparam signed [DEBIT:0]  W_5_x366 =  23'd960;
localparam signed [DEBIT:0]  W_5_x367 =  23'd908;
localparam signed [DEBIT:0]  W_5_x368 =  23'd784;
localparam signed [DEBIT:0]  W_5_x369 =  23'd576;
localparam signed [DEBIT:0]  W_5_x370 =  23'd246;
localparam signed [DEBIT:0]  W_5_x371 = - 23'd3;
localparam signed [DEBIT:0]  W_5_x372 =  23'd76;
localparam signed [DEBIT:0]  W_5_x373 =  23'd279;
localparam signed [DEBIT:0]  W_5_x374 =  23'd204;
localparam signed [DEBIT:0]  W_5_x375 =  23'd132;
localparam signed [DEBIT:0]  W_5_x376 =  23'd255;
localparam signed [DEBIT:0]  W_5_x377 =  23'd293;
localparam signed [DEBIT:0]  W_5_x378 =  23'd86;
localparam signed [DEBIT:0]  W_5_x379 = - 23'd63;
localparam signed [DEBIT:0]  W_5_x380 = - 23'd121;
localparam signed [DEBIT:0]  W_5_x381 = - 23'd293;
localparam signed [DEBIT:0]  W_5_x382 = - 23'd335;
localparam signed [DEBIT:0]  W_5_x383 = - 23'd206;
localparam signed [DEBIT:0]  W_5_x384 = - 23'd77;
localparam signed [DEBIT:0]  W_5_x385 = - 23'd101;
localparam signed [DEBIT:0]  W_5_x386 = - 23'd339;
localparam signed [DEBIT:0]  W_5_x387 = - 23'd625;
localparam signed [DEBIT:0]  W_5_x388 = - 23'd610;
localparam signed [DEBIT:0]  W_5_x389 =  23'd95;
localparam signed [DEBIT:0]  W_5_x390 =  23'd859;
localparam signed [DEBIT:0]  W_5_x391 =  23'd953;
localparam signed [DEBIT:0]  W_5_x392 =  23'd972;
localparam signed [DEBIT:0]  W_5_x393 =  23'd979;
localparam signed [DEBIT:0]  W_5_x394 =  23'd968;
localparam signed [DEBIT:0]  W_5_x395 =  23'd957;
localparam signed [DEBIT:0]  W_5_x396 =  23'd852;
localparam signed [DEBIT:0]  W_5_x397 =  23'd632;
localparam signed [DEBIT:0]  W_5_x398 =  23'd167;
localparam signed [DEBIT:0]  W_5_x399 = - 23'd186;
localparam signed [DEBIT:0]  W_5_x400 = - 23'd129;
localparam signed [DEBIT:0]  W_5_x401 =  23'd121;
localparam signed [DEBIT:0]  W_5_x402 =  23'd190;
localparam signed [DEBIT:0]  W_5_x403 =  23'd241;
localparam signed [DEBIT:0]  W_5_x404 =  23'd120;
localparam signed [DEBIT:0]  W_5_x405 =  23'd168;
localparam signed [DEBIT:0]  W_5_x406 = - 23'd25;
localparam signed [DEBIT:0]  W_5_x407 = - 23'd112;
localparam signed [DEBIT:0]  W_5_x408 = - 23'd104;
localparam signed [DEBIT:0]  W_5_x409 = - 23'd283;
localparam signed [DEBIT:0]  W_5_x410 = - 23'd353;
localparam signed [DEBIT:0]  W_5_x411 = - 23'd249;
localparam signed [DEBIT:0]  W_5_x412 = - 23'd131;
localparam signed [DEBIT:0]  W_5_x413 =  23'd77;
localparam signed [DEBIT:0]  W_5_x414 = - 23'd100;
localparam signed [DEBIT:0]  W_5_x415 = - 23'd297;
localparam signed [DEBIT:0]  W_5_x416 = - 23'd395;
localparam signed [DEBIT:0]  W_5_x417 =  23'd250;
localparam signed [DEBIT:0]  W_5_x418 =  23'd845;
localparam signed [DEBIT:0]  W_5_x419 =  23'd956;
localparam signed [DEBIT:0]  W_5_x420 =  23'd977;
localparam signed [DEBIT:0]  W_5_x421 =  23'd979;
localparam signed [DEBIT:0]  W_5_x422 =  23'd967;
localparam signed [DEBIT:0]  W_5_x423 =  23'd956;
localparam signed [DEBIT:0]  W_5_x424 =  23'd866;
localparam signed [DEBIT:0]  W_5_x425 =  23'd653;
localparam signed [DEBIT:0]  W_5_x426 =  23'd9;
localparam signed [DEBIT:0]  W_5_x427 = - 23'd402;
localparam signed [DEBIT:0]  W_5_x428 = - 23'd412;
localparam signed [DEBIT:0]  W_5_x429 = - 23'd107;
localparam signed [DEBIT:0]  W_5_x430 =  23'd215;
localparam signed [DEBIT:0]  W_5_x431 =  23'd144;
localparam signed [DEBIT:0]  W_5_x432 =  23'd135;
localparam signed [DEBIT:0]  W_5_x433 =  23'd137;
localparam signed [DEBIT:0]  W_5_x434 = - 23'd25;
localparam signed [DEBIT:0]  W_5_x435 = - 23'd106;
localparam signed [DEBIT:0]  W_5_x436 = - 23'd153;
localparam signed [DEBIT:0]  W_5_x437 = - 23'd280;
localparam signed [DEBIT:0]  W_5_x438 = - 23'd271;
localparam signed [DEBIT:0]  W_5_x439 = - 23'd140;
localparam signed [DEBIT:0]  W_5_x440 = - 23'd79;
localparam signed [DEBIT:0]  W_5_x441 = - 23'd62;
localparam signed [DEBIT:0]  W_5_x442 = - 23'd77;
localparam signed [DEBIT:0]  W_5_x443 = - 23'd249;
localparam signed [DEBIT:0]  W_5_x444 = - 23'd201;
localparam signed [DEBIT:0]  W_5_x445 =  23'd333;
localparam signed [DEBIT:0]  W_5_x446 =  23'd811;
localparam signed [DEBIT:0]  W_5_x447 =  23'd939;
localparam signed [DEBIT:0]  W_5_x448 =  23'd979;
localparam signed [DEBIT:0]  W_5_x449 =  23'd980;
localparam signed [DEBIT:0]  W_5_x450 =  23'd962;
localparam signed [DEBIT:0]  W_5_x451 =  23'd955;
localparam signed [DEBIT:0]  W_5_x452 =  23'd880;
localparam signed [DEBIT:0]  W_5_x453 =  23'd664;
localparam signed [DEBIT:0]  W_5_x454 = - 23'd83;
localparam signed [DEBIT:0]  W_5_x455 = - 23'd494;
localparam signed [DEBIT:0]  W_5_x456 = - 23'd501;
localparam signed [DEBIT:0]  W_5_x457 = - 23'd350;
localparam signed [DEBIT:0]  W_5_x458 = - 23'd196;
localparam signed [DEBIT:0]  W_5_x459 = - 23'd129;
localparam signed [DEBIT:0]  W_5_x460 = - 23'd119;
localparam signed [DEBIT:0]  W_5_x461 = - 23'd145;
localparam signed [DEBIT:0]  W_5_x462 = - 23'd166;
localparam signed [DEBIT:0]  W_5_x463 = - 23'd209;
localparam signed [DEBIT:0]  W_5_x464 = - 23'd279;
localparam signed [DEBIT:0]  W_5_x465 = - 23'd319;
localparam signed [DEBIT:0]  W_5_x466 = - 23'd71;
localparam signed [DEBIT:0]  W_5_x467 = - 23'd138;
localparam signed [DEBIT:0]  W_5_x468 = - 23'd92;
localparam signed [DEBIT:0]  W_5_x469 = - 23'd48;
localparam signed [DEBIT:0]  W_5_x470 = - 23'd164;
localparam signed [DEBIT:0]  W_5_x471 = - 23'd202;
localparam signed [DEBIT:0]  W_5_x472 = - 23'd25;
localparam signed [DEBIT:0]  W_5_x473 =  23'd411;
localparam signed [DEBIT:0]  W_5_x474 =  23'd767;
localparam signed [DEBIT:0]  W_5_x475 =  23'd931;
localparam signed [DEBIT:0]  W_5_x476 =  23'd972;
localparam signed [DEBIT:0]  W_5_x477 =  23'd992;
localparam signed [DEBIT:0]  W_5_x478 =  23'd982;
localparam signed [DEBIT:0]  W_5_x479 =  23'd930;
localparam signed [DEBIT:0]  W_5_x480 =  23'd843;
localparam signed [DEBIT:0]  W_5_x481 =  23'd599;
localparam signed [DEBIT:0]  W_5_x482 = - 23'd42;
localparam signed [DEBIT:0]  W_5_x483 = - 23'd63;
localparam signed [DEBIT:0]  W_5_x484 = - 23'd244;
localparam signed [DEBIT:0]  W_5_x485 = - 23'd422;
localparam signed [DEBIT:0]  W_5_x486 = - 23'd488;
localparam signed [DEBIT:0]  W_5_x487 = - 23'd581;
localparam signed [DEBIT:0]  W_5_x488 = - 23'd522;
localparam signed [DEBIT:0]  W_5_x489 = - 23'd391;
localparam signed [DEBIT:0]  W_5_x490 = - 23'd411;
localparam signed [DEBIT:0]  W_5_x491 = - 23'd455;
localparam signed [DEBIT:0]  W_5_x492 = - 23'd320;
localparam signed [DEBIT:0]  W_5_x493 = - 23'd80;
localparam signed [DEBIT:0]  W_5_x494 =  23'd59;
localparam signed [DEBIT:0]  W_5_x495 = - 23'd51;
localparam signed [DEBIT:0]  W_5_x496 = - 23'd117;
localparam signed [DEBIT:0]  W_5_x497 = - 23'd130;
localparam signed [DEBIT:0]  W_5_x498 = - 23'd94;
localparam signed [DEBIT:0]  W_5_x499 = - 23'd165;
localparam signed [DEBIT:0]  W_5_x500 =  23'd110;
localparam signed [DEBIT:0]  W_5_x501 =  23'd452;
localparam signed [DEBIT:0]  W_5_x502 =  23'd775;
localparam signed [DEBIT:0]  W_5_x503 =  23'd929;
localparam signed [DEBIT:0]  W_5_x504 =  23'd980;
localparam signed [DEBIT:0]  W_5_x505 =  23'd976;
localparam signed [DEBIT:0]  W_5_x506 =  23'd976;
localparam signed [DEBIT:0]  W_5_x507 =  23'd934;
localparam signed [DEBIT:0]  W_5_x508 =  23'd797;
localparam signed [DEBIT:0]  W_5_x509 =  23'd514;
localparam signed [DEBIT:0]  W_5_x510 =  23'd27;
localparam signed [DEBIT:0]  W_5_x511 =  23'd247;
localparam signed [DEBIT:0]  W_5_x512 =  23'd93;
localparam signed [DEBIT:0]  W_5_x513 = - 23'd197;
localparam signed [DEBIT:0]  W_5_x514 = - 23'd382;
localparam signed [DEBIT:0]  W_5_x515 = - 23'd549;
localparam signed [DEBIT:0]  W_5_x516 = - 23'd445;
localparam signed [DEBIT:0]  W_5_x517 = - 23'd232;
localparam signed [DEBIT:0]  W_5_x518 = - 23'd171;
localparam signed [DEBIT:0]  W_5_x519 = - 23'd178;
localparam signed [DEBIT:0]  W_5_x520 = - 23'd145;
localparam signed [DEBIT:0]  W_5_x521 = - 23'd22;
localparam signed [DEBIT:0]  W_5_x522 = - 23'd93;
localparam signed [DEBIT:0]  W_5_x523 = - 23'd102;
localparam signed [DEBIT:0]  W_5_x524 = - 23'd106;
localparam signed [DEBIT:0]  W_5_x525 = - 23'd13;
localparam signed [DEBIT:0]  W_5_x526 = - 23'd124;
localparam signed [DEBIT:0]  W_5_x527 = - 23'd150;
localparam signed [DEBIT:0]  W_5_x528 =  23'd142;
localparam signed [DEBIT:0]  W_5_x529 =  23'd494;
localparam signed [DEBIT:0]  W_5_x530 =  23'd808;
localparam signed [DEBIT:0]  W_5_x531 =  23'd940;
localparam signed [DEBIT:0]  W_5_x532 =  23'd988;
localparam signed [DEBIT:0]  W_5_x533 =  23'd989;
localparam signed [DEBIT:0]  W_5_x534 =  23'd968;
localparam signed [DEBIT:0]  W_5_x535 =  23'd911;
localparam signed [DEBIT:0]  W_5_x536 =  23'd702;
localparam signed [DEBIT:0]  W_5_x537 =  23'd413;
localparam signed [DEBIT:0]  W_5_x538 =  23'd61;
localparam signed [DEBIT:0]  W_5_x539 =  23'd206;
localparam signed [DEBIT:0]  W_5_x540 =  23'd225;
localparam signed [DEBIT:0]  W_5_x541 =  23'd90;
localparam signed [DEBIT:0]  W_5_x542 = - 23'd23;
localparam signed [DEBIT:0]  W_5_x543 = - 23'd78;
localparam signed [DEBIT:0]  W_5_x544 =  23'd27;
localparam signed [DEBIT:0]  W_5_x545 =  23'd113;
localparam signed [DEBIT:0]  W_5_x546 =  23'd40;
localparam signed [DEBIT:0]  W_5_x547 = - 23'd12;
localparam signed [DEBIT:0]  W_5_x548 = - 23'd63;
localparam signed [DEBIT:0]  W_5_x549 = - 23'd179;
localparam signed [DEBIT:0]  W_5_x550 = - 23'd205;
localparam signed [DEBIT:0]  W_5_x551 = - 23'd169;
localparam signed [DEBIT:0]  W_5_x552 = - 23'd140;
localparam signed [DEBIT:0]  W_5_x553 = - 23'd133;
localparam signed [DEBIT:0]  W_5_x554 = - 23'd226;
localparam signed [DEBIT:0]  W_5_x555 = - 23'd167;
localparam signed [DEBIT:0]  W_5_x556 =  23'd150;
localparam signed [DEBIT:0]  W_5_x557 =  23'd585;
localparam signed [DEBIT:0]  W_5_x558 =  23'd816;
localparam signed [DEBIT:0]  W_5_x559 =  23'd937;
localparam signed [DEBIT:0]  W_5_x560 =  23'd979;
localparam signed [DEBIT:0]  W_5_x561 =  23'd991;
localparam signed [DEBIT:0]  W_5_x562 =  23'd975;
localparam signed [DEBIT:0]  W_5_x563 =  23'd881;
localparam signed [DEBIT:0]  W_5_x564 =  23'd606;
localparam signed [DEBIT:0]  W_5_x565 =  23'd327;
localparam signed [DEBIT:0]  W_5_x566 =  23'd83;
localparam signed [DEBIT:0]  W_5_x567 =  23'd77;
localparam signed [DEBIT:0]  W_5_x568 =  23'd176;
localparam signed [DEBIT:0]  W_5_x569 =  23'd218;
localparam signed [DEBIT:0]  W_5_x570 =  23'd258;
localparam signed [DEBIT:0]  W_5_x571 =  23'd242;
localparam signed [DEBIT:0]  W_5_x572 =  23'd263;
localparam signed [DEBIT:0]  W_5_x573 =  23'd48;
localparam signed [DEBIT:0]  W_5_x574 = - 23'd27;
localparam signed [DEBIT:0]  W_5_x575 = - 23'd221;
localparam signed [DEBIT:0]  W_5_x576 = - 23'd196;
localparam signed [DEBIT:0]  W_5_x577 = - 23'd109;
localparam signed [DEBIT:0]  W_5_x578 = - 23'd141;
localparam signed [DEBIT:0]  W_5_x579 = - 23'd140;
localparam signed [DEBIT:0]  W_5_x580 = - 23'd67;
localparam signed [DEBIT:0]  W_5_x581 = - 23'd181;
localparam signed [DEBIT:0]  W_5_x582 = - 23'd204;
localparam signed [DEBIT:0]  W_5_x583 = - 23'd96;
localparam signed [DEBIT:0]  W_5_x584 =  23'd263;
localparam signed [DEBIT:0]  W_5_x585 =  23'd639;
localparam signed [DEBIT:0]  W_5_x586 =  23'd850;
localparam signed [DEBIT:0]  W_5_x587 =  23'd960;
localparam signed [DEBIT:0]  W_5_x588 =  23'd976;
localparam signed [DEBIT:0]  W_5_x589 =  23'd979;
localparam signed [DEBIT:0]  W_5_x590 =  23'd973;
localparam signed [DEBIT:0]  W_5_x591 =  23'd885;
localparam signed [DEBIT:0]  W_5_x592 =  23'd653;
localparam signed [DEBIT:0]  W_5_x593 =  23'd306;
localparam signed [DEBIT:0]  W_5_x594 =  23'd13;
localparam signed [DEBIT:0]  W_5_x595 = - 23'd101;
localparam signed [DEBIT:0]  W_5_x596 = - 23'd30;
localparam signed [DEBIT:0]  W_5_x597 =  23'd166;
localparam signed [DEBIT:0]  W_5_x598 =  23'd183;
localparam signed [DEBIT:0]  W_5_x599 =  23'd175;
localparam signed [DEBIT:0]  W_5_x600 =  23'd229;
localparam signed [DEBIT:0]  W_5_x601 =  23'd33;
localparam signed [DEBIT:0]  W_5_x602 = - 23'd4;
localparam signed [DEBIT:0]  W_5_x603 = - 23'd44;
localparam signed [DEBIT:0]  W_5_x604 = - 23'd63;
localparam signed [DEBIT:0]  W_5_x605 = - 23'd40;
localparam signed [DEBIT:0]  W_5_x606 = - 23'd65;
localparam signed [DEBIT:0]  W_5_x607 = - 23'd50;
localparam signed [DEBIT:0]  W_5_x608 = - 23'd4;
localparam signed [DEBIT:0]  W_5_x609 = - 23'd56;
localparam signed [DEBIT:0]  W_5_x610 = - 23'd63;
localparam signed [DEBIT:0]  W_5_x611 =  23'd115;
localparam signed [DEBIT:0]  W_5_x612 =  23'd528;
localparam signed [DEBIT:0]  W_5_x613 =  23'd756;
localparam signed [DEBIT:0]  W_5_x614 =  23'd912;
localparam signed [DEBIT:0]  W_5_x615 =  23'd947;
localparam signed [DEBIT:0]  W_5_x616 =  23'd986;
localparam signed [DEBIT:0]  W_5_x617 =  23'd985;
localparam signed [DEBIT:0]  W_5_x618 =  23'd980;
localparam signed [DEBIT:0]  W_5_x619 =  23'd910;
localparam signed [DEBIT:0]  W_5_x620 =  23'd730;
localparam signed [DEBIT:0]  W_5_x621 =  23'd451;
localparam signed [DEBIT:0]  W_5_x622 =  23'd91;
localparam signed [DEBIT:0]  W_5_x623 = - 23'd191;
localparam signed [DEBIT:0]  W_5_x624 = - 23'd229;
localparam signed [DEBIT:0]  W_5_x625 = - 23'd1;
localparam signed [DEBIT:0]  W_5_x626 =  23'd171;
localparam signed [DEBIT:0]  W_5_x627 =  23'd117;
localparam signed [DEBIT:0]  W_5_x628 =  23'd260;
localparam signed [DEBIT:0]  W_5_x629 =  23'd311;
localparam signed [DEBIT:0]  W_5_x630 =  23'd195;
localparam signed [DEBIT:0]  W_5_x631 =  23'd151;
localparam signed [DEBIT:0]  W_5_x632 =  23'd155;
localparam signed [DEBIT:0]  W_5_x633 =  23'd156;
localparam signed [DEBIT:0]  W_5_x634 =  23'd65;
localparam signed [DEBIT:0]  W_5_x635 =  23'd89;
localparam signed [DEBIT:0]  W_5_x636 =  23'd22;
localparam signed [DEBIT:0]  W_5_x637 = - 23'd74;
localparam signed [DEBIT:0]  W_5_x638 =  23'd61;
localparam signed [DEBIT:0]  W_5_x639 =  23'd418;
localparam signed [DEBIT:0]  W_5_x640 =  23'd721;
localparam signed [DEBIT:0]  W_5_x641 =  23'd869;
localparam signed [DEBIT:0]  W_5_x642 =  23'd947;
localparam signed [DEBIT:0]  W_5_x643 =  23'd972;
localparam signed [DEBIT:0]  W_5_x644 =  23'd984;
localparam signed [DEBIT:0]  W_5_x645 =  23'd984;
localparam signed [DEBIT:0]  W_5_x646 =  23'd973;
localparam signed [DEBIT:0]  W_5_x647 =  23'd953;
localparam signed [DEBIT:0]  W_5_x648 =  23'd872;
localparam signed [DEBIT:0]  W_5_x649 =  23'd699;
localparam signed [DEBIT:0]  W_5_x650 =  23'd427;
localparam signed [DEBIT:0]  W_5_x651 =  23'd122;
localparam signed [DEBIT:0]  W_5_x652 = - 23'd109;
localparam signed [DEBIT:0]  W_5_x653 = - 23'd70;
localparam signed [DEBIT:0]  W_5_x654 =  23'd28;
localparam signed [DEBIT:0]  W_5_x655 =  23'd62;
localparam signed [DEBIT:0]  W_5_x656 =  23'd141;
localparam signed [DEBIT:0]  W_5_x657 =  23'd198;
localparam signed [DEBIT:0]  W_5_x658 =  23'd127;
localparam signed [DEBIT:0]  W_5_x659 =  23'd164;
localparam signed [DEBIT:0]  W_5_x660 =  23'd177;
localparam signed [DEBIT:0]  W_5_x661 =  23'd195;
localparam signed [DEBIT:0]  W_5_x662 =  23'd74;
localparam signed [DEBIT:0]  W_5_x663 = - 23'd88;
localparam signed [DEBIT:0]  W_5_x664 = - 23'd32;
localparam signed [DEBIT:0]  W_5_x665 =  23'd117;
localparam signed [DEBIT:0]  W_5_x666 =  23'd403;
localparam signed [DEBIT:0]  W_5_x667 =  23'd687;
localparam signed [DEBIT:0]  W_5_x668 =  23'd847;
localparam signed [DEBIT:0]  W_5_x669 =  23'd931;
localparam signed [DEBIT:0]  W_5_x670 =  23'd968;
localparam signed [DEBIT:0]  W_5_x671 =  23'd978;
localparam signed [DEBIT:0]  W_5_x672 =  23'd973;
localparam signed [DEBIT:0]  W_5_x673 =  23'd980;
localparam signed [DEBIT:0]  W_5_x674 =  23'd966;
localparam signed [DEBIT:0]  W_5_x675 =  23'd960;
localparam signed [DEBIT:0]  W_5_x676 =  23'd940;
localparam signed [DEBIT:0]  W_5_x677 =  23'd869;
localparam signed [DEBIT:0]  W_5_x678 =  23'd725;
localparam signed [DEBIT:0]  W_5_x679 =  23'd519;
localparam signed [DEBIT:0]  W_5_x680 =  23'd301;
localparam signed [DEBIT:0]  W_5_x681 =  23'd151;
localparam signed [DEBIT:0]  W_5_x682 =  23'd40;
localparam signed [DEBIT:0]  W_5_x683 =  23'd37;
localparam signed [DEBIT:0]  W_5_x684 =  23'd105;
localparam signed [DEBIT:0]  W_5_x685 =  23'd165;
localparam signed [DEBIT:0]  W_5_x686 =  23'd117;
localparam signed [DEBIT:0]  W_5_x687 =  23'd109;
localparam signed [DEBIT:0]  W_5_x688 =  23'd72;
localparam signed [DEBIT:0]  W_5_x689 =  23'd15;
localparam signed [DEBIT:0]  W_5_x690 =  23'd22;
localparam signed [DEBIT:0]  W_5_x691 =  23'd106;
localparam signed [DEBIT:0]  W_5_x692 =  23'd300;
localparam signed [DEBIT:0]  W_5_x693 =  23'd461;
localparam signed [DEBIT:0]  W_5_x694 =  23'd652;
localparam signed [DEBIT:0]  W_5_x695 =  23'd835;
localparam signed [DEBIT:0]  W_5_x696 =  23'd907;
localparam signed [DEBIT:0]  W_5_x697 =  23'd953;
localparam signed [DEBIT:0]  W_5_x698 =  23'd985;
localparam signed [DEBIT:0]  W_5_x699 =  23'd982;
localparam signed [DEBIT:0]  W_5_x700 =  23'd980;
localparam signed [DEBIT:0]  W_5_x701 =  23'd971;
localparam signed [DEBIT:0]  W_5_x702 =  23'd974;
localparam signed [DEBIT:0]  W_5_x703 =  23'd979;
localparam signed [DEBIT:0]  W_5_x704 =  23'd972;
localparam signed [DEBIT:0]  W_5_x705 =  23'd943;
localparam signed [DEBIT:0]  W_5_x706 =  23'd907;
localparam signed [DEBIT:0]  W_5_x707 =  23'd820;
localparam signed [DEBIT:0]  W_5_x708 =  23'd727;
localparam signed [DEBIT:0]  W_5_x709 =  23'd615;
localparam signed [DEBIT:0]  W_5_x710 =  23'd500;
localparam signed [DEBIT:0]  W_5_x711 =  23'd412;
localparam signed [DEBIT:0]  W_5_x712 =  23'd411;
localparam signed [DEBIT:0]  W_5_x713 =  23'd353;
localparam signed [DEBIT:0]  W_5_x714 =  23'd278;
localparam signed [DEBIT:0]  W_5_x715 =  23'd242;
localparam signed [DEBIT:0]  W_5_x716 =  23'd296;
localparam signed [DEBIT:0]  W_5_x717 =  23'd289;
localparam signed [DEBIT:0]  W_5_x718 =  23'd341;
localparam signed [DEBIT:0]  W_5_x719 =  23'd426;
localparam signed [DEBIT:0]  W_5_x720 =  23'd577;
localparam signed [DEBIT:0]  W_5_x721 =  23'd697;
localparam signed [DEBIT:0]  W_5_x722 =  23'd814;
localparam signed [DEBIT:0]  W_5_x723 =  23'd892;
localparam signed [DEBIT:0]  W_5_x724 =  23'd943;
localparam signed [DEBIT:0]  W_5_x725 =  23'd983;
localparam signed [DEBIT:0]  W_5_x726 =  23'd973;
localparam signed [DEBIT:0]  W_5_x727 =  23'd993;
localparam signed [DEBIT:0]  W_5_x728 =  23'd978;
localparam signed [DEBIT:0]  W_5_x729 =  23'd974;
localparam signed [DEBIT:0]  W_5_x730 =  23'd978;
localparam signed [DEBIT:0]  W_5_x731 =  23'd976;
localparam signed [DEBIT:0]  W_5_x732 =  23'd987;
localparam signed [DEBIT:0]  W_5_x733 =  23'd970;
localparam signed [DEBIT:0]  W_5_x734 =  23'd955;
localparam signed [DEBIT:0]  W_5_x735 =  23'd901;
localparam signed [DEBIT:0]  W_5_x736 =  23'd879;
localparam signed [DEBIT:0]  W_5_x737 =  23'd834;
localparam signed [DEBIT:0]  W_5_x738 =  23'd788;
localparam signed [DEBIT:0]  W_5_x739 =  23'd772;
localparam signed [DEBIT:0]  W_5_x740 =  23'd749;
localparam signed [DEBIT:0]  W_5_x741 =  23'd710;
localparam signed [DEBIT:0]  W_5_x742 =  23'd643;
localparam signed [DEBIT:0]  W_5_x743 =  23'd599;
localparam signed [DEBIT:0]  W_5_x744 =  23'd605;
localparam signed [DEBIT:0]  W_5_x745 =  23'd589;
localparam signed [DEBIT:0]  W_5_x746 =  23'd589;
localparam signed [DEBIT:0]  W_5_x747 =  23'd626;
localparam signed [DEBIT:0]  W_5_x748 =  23'd743;
localparam signed [DEBIT:0]  W_5_x749 =  23'd862;
localparam signed [DEBIT:0]  W_5_x750 =  23'd897;
localparam signed [DEBIT:0]  W_5_x751 =  23'd941;
localparam signed [DEBIT:0]  W_5_x752 =  23'd976;
localparam signed [DEBIT:0]  W_5_x753 =  23'd988;
localparam signed [DEBIT:0]  W_5_x754 =  23'd979;
localparam signed [DEBIT:0]  W_5_x755 =  23'd973;
localparam signed [DEBIT:0]  W_5_x756 =  23'd974;
localparam signed [DEBIT:0]  W_5_x757 =  23'd978;
localparam signed [DEBIT:0]  W_5_x758 =  23'd973;
localparam signed [DEBIT:0]  W_5_x759 =  23'd968;
localparam signed [DEBIT:0]  W_5_x760 =  23'd978;
localparam signed [DEBIT:0]  W_5_x761 =  23'd982;
localparam signed [DEBIT:0]  W_5_x762 =  23'd968;
localparam signed [DEBIT:0]  W_5_x763 =  23'd960;
localparam signed [DEBIT:0]  W_5_x764 =  23'd957;
localparam signed [DEBIT:0]  W_5_x765 =  23'd964;
localparam signed [DEBIT:0]  W_5_x766 =  23'd976;
localparam signed [DEBIT:0]  W_5_x767 =  23'd970;
localparam signed [DEBIT:0]  W_5_x768 =  23'd940;
localparam signed [DEBIT:0]  W_5_x769 =  23'd897;
localparam signed [DEBIT:0]  W_5_x770 =  23'd878;
localparam signed [DEBIT:0]  W_5_x771 =  23'd853;
localparam signed [DEBIT:0]  W_5_x772 =  23'd856;
localparam signed [DEBIT:0]  W_5_x773 =  23'd853;
localparam signed [DEBIT:0]  W_5_x774 =  23'd845;
localparam signed [DEBIT:0]  W_5_x775 =  23'd847;
localparam signed [DEBIT:0]  W_5_x776 =  23'd897;
localparam signed [DEBIT:0]  W_5_x777 =  23'd930;
localparam signed [DEBIT:0]  W_5_x778 =  23'd953;
localparam signed [DEBIT:0]  W_5_x779 =  23'd966;
localparam signed [DEBIT:0]  W_5_x780 =  23'd976;
localparam signed [DEBIT:0]  W_5_x781 =  23'd975;
localparam signed [DEBIT:0]  W_5_x782 =  23'd978;
localparam signed [DEBIT:0]  W_5_x783 =  23'd986;
localparam signed [DEBIT:0]  W_5_x784 =  23'd981;
localparam signed [DEBIT:0]  W_6_x1 =  23'd968;
localparam signed [DEBIT:0]  W_6_x2 =  23'd968;
localparam signed [DEBIT:0]  W_6_x3 =  23'd970;
localparam signed [DEBIT:0]  W_6_x4 =  23'd968;
localparam signed [DEBIT:0]  W_6_x5 =  23'd968;
localparam signed [DEBIT:0]  W_6_x6 =  23'd961;
localparam signed [DEBIT:0]  W_6_x7 =  23'd971;
localparam signed [DEBIT:0]  W_6_x8 =  23'd972;
localparam signed [DEBIT:0]  W_6_x9 =  23'd971;
localparam signed [DEBIT:0]  W_6_x10 =  23'd956;
localparam signed [DEBIT:0]  W_6_x11 =  23'd968;
localparam signed [DEBIT:0]  W_6_x12 =  23'd962;
localparam signed [DEBIT:0]  W_6_x13 =  23'd972;
localparam signed [DEBIT:0]  W_6_x14 =  23'd974;
localparam signed [DEBIT:0]  W_6_x15 =  23'd963;
localparam signed [DEBIT:0]  W_6_x16 =  23'd969;
localparam signed [DEBIT:0]  W_6_x17 =  23'd969;
localparam signed [DEBIT:0]  W_6_x18 =  23'd977;
localparam signed [DEBIT:0]  W_6_x19 =  23'd970;
localparam signed [DEBIT:0]  W_6_x20 =  23'd979;
localparam signed [DEBIT:0]  W_6_x21 =  23'd960;
localparam signed [DEBIT:0]  W_6_x22 =  23'd964;
localparam signed [DEBIT:0]  W_6_x23 =  23'd978;
localparam signed [DEBIT:0]  W_6_x24 =  23'd977;
localparam signed [DEBIT:0]  W_6_x25 =  23'd962;
localparam signed [DEBIT:0]  W_6_x26 =  23'd961;
localparam signed [DEBIT:0]  W_6_x27 =  23'd980;
localparam signed [DEBIT:0]  W_6_x28 =  23'd970;
localparam signed [DEBIT:0]  W_6_x29 =  23'd974;
localparam signed [DEBIT:0]  W_6_x30 =  23'd973;
localparam signed [DEBIT:0]  W_6_x31 =  23'd965;
localparam signed [DEBIT:0]  W_6_x32 =  23'd962;
localparam signed [DEBIT:0]  W_6_x33 =  23'd976;
localparam signed [DEBIT:0]  W_6_x34 =  23'd968;
localparam signed [DEBIT:0]  W_6_x35 =  23'd965;
localparam signed [DEBIT:0]  W_6_x36 =  23'd972;
localparam signed [DEBIT:0]  W_6_x37 =  23'd979;
localparam signed [DEBIT:0]  W_6_x38 =  23'd963;
localparam signed [DEBIT:0]  W_6_x39 =  23'd960;
localparam signed [DEBIT:0]  W_6_x40 =  23'd956;
localparam signed [DEBIT:0]  W_6_x41 =  23'd958;
localparam signed [DEBIT:0]  W_6_x42 =  23'd967;
localparam signed [DEBIT:0]  W_6_x43 =  23'd965;
localparam signed [DEBIT:0]  W_6_x44 =  23'd961;
localparam signed [DEBIT:0]  W_6_x45 =  23'd947;
localparam signed [DEBIT:0]  W_6_x46 =  23'd967;
localparam signed [DEBIT:0]  W_6_x47 =  23'd965;
localparam signed [DEBIT:0]  W_6_x48 =  23'd968;
localparam signed [DEBIT:0]  W_6_x49 =  23'd977;
localparam signed [DEBIT:0]  W_6_x50 =  23'd972;
localparam signed [DEBIT:0]  W_6_x51 =  23'd967;
localparam signed [DEBIT:0]  W_6_x52 =  23'd975;
localparam signed [DEBIT:0]  W_6_x53 =  23'd976;
localparam signed [DEBIT:0]  W_6_x54 =  23'd975;
localparam signed [DEBIT:0]  W_6_x55 =  23'd978;
localparam signed [DEBIT:0]  W_6_x56 =  23'd976;
localparam signed [DEBIT:0]  W_6_x57 =  23'd968;
localparam signed [DEBIT:0]  W_6_x58 =  23'd962;
localparam signed [DEBIT:0]  W_6_x59 =  23'd973;
localparam signed [DEBIT:0]  W_6_x60 =  23'd967;
localparam signed [DEBIT:0]  W_6_x61 =  23'd974;
localparam signed [DEBIT:0]  W_6_x62 =  23'd974;
localparam signed [DEBIT:0]  W_6_x63 =  23'd964;
localparam signed [DEBIT:0]  W_6_x64 =  23'd951;
localparam signed [DEBIT:0]  W_6_x65 =  23'd948;
localparam signed [DEBIT:0]  W_6_x66 =  23'd917;
localparam signed [DEBIT:0]  W_6_x67 =  23'd931;
localparam signed [DEBIT:0]  W_6_x68 =  23'd909;
localparam signed [DEBIT:0]  W_6_x69 =  23'd849;
localparam signed [DEBIT:0]  W_6_x70 =  23'd838;
localparam signed [DEBIT:0]  W_6_x71 =  23'd822;
localparam signed [DEBIT:0]  W_6_x72 =  23'd796;
localparam signed [DEBIT:0]  W_6_x73 =  23'd851;
localparam signed [DEBIT:0]  W_6_x74 =  23'd938;
localparam signed [DEBIT:0]  W_6_x75 =  23'd1021;
localparam signed [DEBIT:0]  W_6_x76 =  23'd1044;
localparam signed [DEBIT:0]  W_6_x77 =  23'd1013;
localparam signed [DEBIT:0]  W_6_x78 =  23'd1017;
localparam signed [DEBIT:0]  W_6_x79 =  23'd993;
localparam signed [DEBIT:0]  W_6_x80 =  23'd980;
localparam signed [DEBIT:0]  W_6_x81 =  23'd967;
localparam signed [DEBIT:0]  W_6_x82 =  23'd963;
localparam signed [DEBIT:0]  W_6_x83 =  23'd968;
localparam signed [DEBIT:0]  W_6_x84 =  23'd973;
localparam signed [DEBIT:0]  W_6_x85 =  23'd968;
localparam signed [DEBIT:0]  W_6_x86 =  23'd975;
localparam signed [DEBIT:0]  W_6_x87 =  23'd972;
localparam signed [DEBIT:0]  W_6_x88 =  23'd970;
localparam signed [DEBIT:0]  W_6_x89 =  23'd974;
localparam signed [DEBIT:0]  W_6_x90 =  23'd955;
localparam signed [DEBIT:0]  W_6_x91 =  23'd896;
localparam signed [DEBIT:0]  W_6_x92 =  23'd791;
localparam signed [DEBIT:0]  W_6_x93 =  23'd682;
localparam signed [DEBIT:0]  W_6_x94 =  23'd597;
localparam signed [DEBIT:0]  W_6_x95 =  23'd544;
localparam signed [DEBIT:0]  W_6_x96 =  23'd445;
localparam signed [DEBIT:0]  W_6_x97 =  23'd350;
localparam signed [DEBIT:0]  W_6_x98 =  23'd414;
localparam signed [DEBIT:0]  W_6_x99 =  23'd464;
localparam signed [DEBIT:0]  W_6_x100 =  23'd522;
localparam signed [DEBIT:0]  W_6_x101 =  23'd657;
localparam signed [DEBIT:0]  W_6_x102 =  23'd768;
localparam signed [DEBIT:0]  W_6_x103 =  23'd906;
localparam signed [DEBIT:0]  W_6_x104 =  23'd1018;
localparam signed [DEBIT:0]  W_6_x105 =  23'd1035;
localparam signed [DEBIT:0]  W_6_x106 =  23'd1002;
localparam signed [DEBIT:0]  W_6_x107 =  23'd943;
localparam signed [DEBIT:0]  W_6_x108 =  23'd952;
localparam signed [DEBIT:0]  W_6_x109 =  23'd987;
localparam signed [DEBIT:0]  W_6_x110 =  23'd974;
localparam signed [DEBIT:0]  W_6_x111 =  23'd965;
localparam signed [DEBIT:0]  W_6_x112 =  23'd969;
localparam signed [DEBIT:0]  W_6_x113 =  23'd974;
localparam signed [DEBIT:0]  W_6_x114 =  23'd965;
localparam signed [DEBIT:0]  W_6_x115 =  23'd969;
localparam signed [DEBIT:0]  W_6_x116 =  23'd973;
localparam signed [DEBIT:0]  W_6_x117 =  23'd967;
localparam signed [DEBIT:0]  W_6_x118 =  23'd881;
localparam signed [DEBIT:0]  W_6_x119 =  23'd736;
localparam signed [DEBIT:0]  W_6_x120 =  23'd518;
localparam signed [DEBIT:0]  W_6_x121 =  23'd315;
localparam signed [DEBIT:0]  W_6_x122 =  23'd179;
localparam signed [DEBIT:0]  W_6_x123 =  23'd120;
localparam signed [DEBIT:0]  W_6_x124 = - 23'd12;
localparam signed [DEBIT:0]  W_6_x125 = - 23'd79;
localparam signed [DEBIT:0]  W_6_x126 = - 23'd6;
localparam signed [DEBIT:0]  W_6_x127 =  23'd105;
localparam signed [DEBIT:0]  W_6_x128 =  23'd116;
localparam signed [DEBIT:0]  W_6_x129 =  23'd120;
localparam signed [DEBIT:0]  W_6_x130 =  23'd343;
localparam signed [DEBIT:0]  W_6_x131 =  23'd478;
localparam signed [DEBIT:0]  W_6_x132 =  23'd558;
localparam signed [DEBIT:0]  W_6_x133 =  23'd627;
localparam signed [DEBIT:0]  W_6_x134 =  23'd638;
localparam signed [DEBIT:0]  W_6_x135 =  23'd678;
localparam signed [DEBIT:0]  W_6_x136 =  23'd816;
localparam signed [DEBIT:0]  W_6_x137 =  23'd897;
localparam signed [DEBIT:0]  W_6_x138 =  23'd944;
localparam signed [DEBIT:0]  W_6_x139 =  23'd959;
localparam signed [DEBIT:0]  W_6_x140 =  23'd963;
localparam signed [DEBIT:0]  W_6_x141 =  23'd970;
localparam signed [DEBIT:0]  W_6_x142 =  23'd975;
localparam signed [DEBIT:0]  W_6_x143 =  23'd975;
localparam signed [DEBIT:0]  W_6_x144 =  23'd961;
localparam signed [DEBIT:0]  W_6_x145 =  23'd908;
localparam signed [DEBIT:0]  W_6_x146 =  23'd726;
localparam signed [DEBIT:0]  W_6_x147 =  23'd416;
localparam signed [DEBIT:0]  W_6_x148 =  23'd125;
localparam signed [DEBIT:0]  W_6_x149 = - 23'd38;
localparam signed [DEBIT:0]  W_6_x150 = - 23'd52;
localparam signed [DEBIT:0]  W_6_x151 = - 23'd84;
localparam signed [DEBIT:0]  W_6_x152 = - 23'd211;
localparam signed [DEBIT:0]  W_6_x153 = - 23'd165;
localparam signed [DEBIT:0]  W_6_x154 = - 23'd281;
localparam signed [DEBIT:0]  W_6_x155 = - 23'd54;
localparam signed [DEBIT:0]  W_6_x156 = - 23'd82;
localparam signed [DEBIT:0]  W_6_x157 = - 23'd95;
localparam signed [DEBIT:0]  W_6_x158 = - 23'd61;
localparam signed [DEBIT:0]  W_6_x159 =  23'd52;
localparam signed [DEBIT:0]  W_6_x160 =  23'd95;
localparam signed [DEBIT:0]  W_6_x161 =  23'd71;
localparam signed [DEBIT:0]  W_6_x162 =  23'd59;
localparam signed [DEBIT:0]  W_6_x163 =  23'd293;
localparam signed [DEBIT:0]  W_6_x164 =  23'd578;
localparam signed [DEBIT:0]  W_6_x165 =  23'd768;
localparam signed [DEBIT:0]  W_6_x166 =  23'd853;
localparam signed [DEBIT:0]  W_6_x167 =  23'd959;
localparam signed [DEBIT:0]  W_6_x168 =  23'd965;
localparam signed [DEBIT:0]  W_6_x169 =  23'd977;
localparam signed [DEBIT:0]  W_6_x170 =  23'd962;
localparam signed [DEBIT:0]  W_6_x171 =  23'd958;
localparam signed [DEBIT:0]  W_6_x172 =  23'd922;
localparam signed [DEBIT:0]  W_6_x173 =  23'd807;
localparam signed [DEBIT:0]  W_6_x174 =  23'd521;
localparam signed [DEBIT:0]  W_6_x175 =  23'd190;
localparam signed [DEBIT:0]  W_6_x176 = - 23'd63;
localparam signed [DEBIT:0]  W_6_x177 = - 23'd149;
localparam signed [DEBIT:0]  W_6_x178 = - 23'd124;
localparam signed [DEBIT:0]  W_6_x179 = - 23'd207;
localparam signed [DEBIT:0]  W_6_x180 = - 23'd148;
localparam signed [DEBIT:0]  W_6_x181 = - 23'd156;
localparam signed [DEBIT:0]  W_6_x182 = - 23'd165;
localparam signed [DEBIT:0]  W_6_x183 = - 23'd134;
localparam signed [DEBIT:0]  W_6_x184 = - 23'd142;
localparam signed [DEBIT:0]  W_6_x185 = - 23'd79;
localparam signed [DEBIT:0]  W_6_x186 = - 23'd117;
localparam signed [DEBIT:0]  W_6_x187 = - 23'd189;
localparam signed [DEBIT:0]  W_6_x188 = - 23'd208;
localparam signed [DEBIT:0]  W_6_x189 = - 23'd369;
localparam signed [DEBIT:0]  W_6_x190 = - 23'd342;
localparam signed [DEBIT:0]  W_6_x191 = - 23'd82;
localparam signed [DEBIT:0]  W_6_x192 =  23'd283;
localparam signed [DEBIT:0]  W_6_x193 =  23'd542;
localparam signed [DEBIT:0]  W_6_x194 =  23'd746;
localparam signed [DEBIT:0]  W_6_x195 =  23'd907;
localparam signed [DEBIT:0]  W_6_x196 =  23'd965;
localparam signed [DEBIT:0]  W_6_x197 =  23'd975;
localparam signed [DEBIT:0]  W_6_x198 =  23'd970;
localparam signed [DEBIT:0]  W_6_x199 =  23'd940;
localparam signed [DEBIT:0]  W_6_x200 =  23'd820;
localparam signed [DEBIT:0]  W_6_x201 =  23'd628;
localparam signed [DEBIT:0]  W_6_x202 =  23'd319;
localparam signed [DEBIT:0]  W_6_x203 =  23'd34;
localparam signed [DEBIT:0]  W_6_x204 = - 23'd110;
localparam signed [DEBIT:0]  W_6_x205 = - 23'd94;
localparam signed [DEBIT:0]  W_6_x206 = - 23'd104;
localparam signed [DEBIT:0]  W_6_x207 = - 23'd5;
localparam signed [DEBIT:0]  W_6_x208 = - 23'd47;
localparam signed [DEBIT:0]  W_6_x209 = - 23'd127;
localparam signed [DEBIT:0]  W_6_x210 = - 23'd222;
localparam signed [DEBIT:0]  W_6_x211 = - 23'd255;
localparam signed [DEBIT:0]  W_6_x212 = - 23'd274;
localparam signed [DEBIT:0]  W_6_x213 = - 23'd277;
localparam signed [DEBIT:0]  W_6_x214 = - 23'd261;
localparam signed [DEBIT:0]  W_6_x215 = - 23'd290;
localparam signed [DEBIT:0]  W_6_x216 = - 23'd323;
localparam signed [DEBIT:0]  W_6_x217 = - 23'd493;
localparam signed [DEBIT:0]  W_6_x218 = - 23'd503;
localparam signed [DEBIT:0]  W_6_x219 = - 23'd364;
localparam signed [DEBIT:0]  W_6_x220 =  23'd5;
localparam signed [DEBIT:0]  W_6_x221 =  23'd420;
localparam signed [DEBIT:0]  W_6_x222 =  23'd705;
localparam signed [DEBIT:0]  W_6_x223 =  23'd882;
localparam signed [DEBIT:0]  W_6_x224 =  23'd965;
localparam signed [DEBIT:0]  W_6_x225 =  23'd974;
localparam signed [DEBIT:0]  W_6_x226 =  23'd940;
localparam signed [DEBIT:0]  W_6_x227 =  23'd857;
localparam signed [DEBIT:0]  W_6_x228 =  23'd691;
localparam signed [DEBIT:0]  W_6_x229 =  23'd385;
localparam signed [DEBIT:0]  W_6_x230 =  23'd113;
localparam signed [DEBIT:0]  W_6_x231 = - 23'd124;
localparam signed [DEBIT:0]  W_6_x232 = - 23'd197;
localparam signed [DEBIT:0]  W_6_x233 = - 23'd188;
localparam signed [DEBIT:0]  W_6_x234 = - 23'd63;
localparam signed [DEBIT:0]  W_6_x235 = - 23'd85;
localparam signed [DEBIT:0]  W_6_x236 = - 23'd118;
localparam signed [DEBIT:0]  W_6_x237 = - 23'd181;
localparam signed [DEBIT:0]  W_6_x238 = - 23'd296;
localparam signed [DEBIT:0]  W_6_x239 = - 23'd327;
localparam signed [DEBIT:0]  W_6_x240 = - 23'd329;
localparam signed [DEBIT:0]  W_6_x241 = - 23'd346;
localparam signed [DEBIT:0]  W_6_x242 = - 23'd428;
localparam signed [DEBIT:0]  W_6_x243 = - 23'd536;
localparam signed [DEBIT:0]  W_6_x244 = - 23'd541;
localparam signed [DEBIT:0]  W_6_x245 = - 23'd570;
localparam signed [DEBIT:0]  W_6_x246 = - 23'd660;
localparam signed [DEBIT:0]  W_6_x247 = - 23'd550;
localparam signed [DEBIT:0]  W_6_x248 = - 23'd140;
localparam signed [DEBIT:0]  W_6_x249 =  23'd362;
localparam signed [DEBIT:0]  W_6_x250 =  23'd694;
localparam signed [DEBIT:0]  W_6_x251 =  23'd859;
localparam signed [DEBIT:0]  W_6_x252 =  23'd964;
localparam signed [DEBIT:0]  W_6_x253 =  23'd970;
localparam signed [DEBIT:0]  W_6_x254 =  23'd922;
localparam signed [DEBIT:0]  W_6_x255 =  23'd827;
localparam signed [DEBIT:0]  W_6_x256 =  23'd612;
localparam signed [DEBIT:0]  W_6_x257 =  23'd332;
localparam signed [DEBIT:0]  W_6_x258 =  23'd6;
localparam signed [DEBIT:0]  W_6_x259 = - 23'd240;
localparam signed [DEBIT:0]  W_6_x260 = - 23'd244;
localparam signed [DEBIT:0]  W_6_x261 = - 23'd160;
localparam signed [DEBIT:0]  W_6_x262 = - 23'd137;
localparam signed [DEBIT:0]  W_6_x263 = - 23'd143;
localparam signed [DEBIT:0]  W_6_x264 = - 23'd127;
localparam signed [DEBIT:0]  W_6_x265 = - 23'd159;
localparam signed [DEBIT:0]  W_6_x266 = - 23'd267;
localparam signed [DEBIT:0]  W_6_x267 = - 23'd332;
localparam signed [DEBIT:0]  W_6_x268 = - 23'd285;
localparam signed [DEBIT:0]  W_6_x269 = - 23'd460;
localparam signed [DEBIT:0]  W_6_x270 = - 23'd584;
localparam signed [DEBIT:0]  W_6_x271 = - 23'd607;
localparam signed [DEBIT:0]  W_6_x272 = - 23'd483;
localparam signed [DEBIT:0]  W_6_x273 = - 23'd473;
localparam signed [DEBIT:0]  W_6_x274 = - 23'd568;
localparam signed [DEBIT:0]  W_6_x275 = - 23'd527;
localparam signed [DEBIT:0]  W_6_x276 = - 23'd141;
localparam signed [DEBIT:0]  W_6_x277 =  23'd357;
localparam signed [DEBIT:0]  W_6_x278 =  23'd695;
localparam signed [DEBIT:0]  W_6_x279 =  23'd864;
localparam signed [DEBIT:0]  W_6_x280 =  23'd959;
localparam signed [DEBIT:0]  W_6_x281 =  23'd978;
localparam signed [DEBIT:0]  W_6_x282 =  23'd909;
localparam signed [DEBIT:0]  W_6_x283 =  23'd841;
localparam signed [DEBIT:0]  W_6_x284 =  23'd631;
localparam signed [DEBIT:0]  W_6_x285 =  23'd343;
localparam signed [DEBIT:0]  W_6_x286 =  23'd27;
localparam signed [DEBIT:0]  W_6_x287 = - 23'd229;
localparam signed [DEBIT:0]  W_6_x288 = - 23'd183;
localparam signed [DEBIT:0]  W_6_x289 = - 23'd42;
localparam signed [DEBIT:0]  W_6_x290 = - 23'd26;
localparam signed [DEBIT:0]  W_6_x291 = - 23'd167;
localparam signed [DEBIT:0]  W_6_x292 = - 23'd113;
localparam signed [DEBIT:0]  W_6_x293 = - 23'd94;
localparam signed [DEBIT:0]  W_6_x294 = - 23'd100;
localparam signed [DEBIT:0]  W_6_x295 = - 23'd255;
localparam signed [DEBIT:0]  W_6_x296 = - 23'd401;
localparam signed [DEBIT:0]  W_6_x297 = - 23'd584;
localparam signed [DEBIT:0]  W_6_x298 = - 23'd465;
localparam signed [DEBIT:0]  W_6_x299 = - 23'd416;
localparam signed [DEBIT:0]  W_6_x300 = - 23'd385;
localparam signed [DEBIT:0]  W_6_x301 = - 23'd368;
localparam signed [DEBIT:0]  W_6_x302 = - 23'd384;
localparam signed [DEBIT:0]  W_6_x303 = - 23'd351;
localparam signed [DEBIT:0]  W_6_x304 = - 23'd3;
localparam signed [DEBIT:0]  W_6_x305 =  23'd438;
localparam signed [DEBIT:0]  W_6_x306 =  23'd740;
localparam signed [DEBIT:0]  W_6_x307 =  23'd880;
localparam signed [DEBIT:0]  W_6_x308 =  23'd945;
localparam signed [DEBIT:0]  W_6_x309 =  23'd967;
localparam signed [DEBIT:0]  W_6_x310 =  23'd929;
localparam signed [DEBIT:0]  W_6_x311 =  23'd851;
localparam signed [DEBIT:0]  W_6_x312 =  23'd664;
localparam signed [DEBIT:0]  W_6_x313 =  23'd404;
localparam signed [DEBIT:0]  W_6_x314 =  23'd65;
localparam signed [DEBIT:0]  W_6_x315 = - 23'd173;
localparam signed [DEBIT:0]  W_6_x316 = - 23'd122;
localparam signed [DEBIT:0]  W_6_x317 =  23'd119;
localparam signed [DEBIT:0]  W_6_x318 =  23'd23;
localparam signed [DEBIT:0]  W_6_x319 = - 23'd94;
localparam signed [DEBIT:0]  W_6_x320 = - 23'd41;
localparam signed [DEBIT:0]  W_6_x321 =  23'd59;
localparam signed [DEBIT:0]  W_6_x322 =  23'd20;
localparam signed [DEBIT:0]  W_6_x323 = - 23'd274;
localparam signed [DEBIT:0]  W_6_x324 = - 23'd413;
localparam signed [DEBIT:0]  W_6_x325 = - 23'd318;
localparam signed [DEBIT:0]  W_6_x326 = - 23'd163;
localparam signed [DEBIT:0]  W_6_x327 = - 23'd91;
localparam signed [DEBIT:0]  W_6_x328 = - 23'd210;
localparam signed [DEBIT:0]  W_6_x329 = - 23'd320;
localparam signed [DEBIT:0]  W_6_x330 = - 23'd138;
localparam signed [DEBIT:0]  W_6_x331 = - 23'd90;
localparam signed [DEBIT:0]  W_6_x332 =  23'd209;
localparam signed [DEBIT:0]  W_6_x333 =  23'd528;
localparam signed [DEBIT:0]  W_6_x334 =  23'd792;
localparam signed [DEBIT:0]  W_6_x335 =  23'd899;
localparam signed [DEBIT:0]  W_6_x336 =  23'd955;
localparam signed [DEBIT:0]  W_6_x337 =  23'd966;
localparam signed [DEBIT:0]  W_6_x338 =  23'd942;
localparam signed [DEBIT:0]  W_6_x339 =  23'd875;
localparam signed [DEBIT:0]  W_6_x340 =  23'd736;
localparam signed [DEBIT:0]  W_6_x341 =  23'd432;
localparam signed [DEBIT:0]  W_6_x342 =  23'd30;
localparam signed [DEBIT:0]  W_6_x343 = - 23'd142;
localparam signed [DEBIT:0]  W_6_x344 =  23'd33;
localparam signed [DEBIT:0]  W_6_x345 =  23'd218;
localparam signed [DEBIT:0]  W_6_x346 =  23'd107;
localparam signed [DEBIT:0]  W_6_x347 = - 23'd22;
localparam signed [DEBIT:0]  W_6_x348 =  23'd104;
localparam signed [DEBIT:0]  W_6_x349 =  23'd301;
localparam signed [DEBIT:0]  W_6_x350 =  23'd112;
localparam signed [DEBIT:0]  W_6_x351 = - 23'd262;
localparam signed [DEBIT:0]  W_6_x352 = - 23'd232;
localparam signed [DEBIT:0]  W_6_x353 = - 23'd29;
localparam signed [DEBIT:0]  W_6_x354 =  23'd78;
localparam signed [DEBIT:0]  W_6_x355 = - 23'd3;
localparam signed [DEBIT:0]  W_6_x356 = - 23'd177;
localparam signed [DEBIT:0]  W_6_x357 = - 23'd150;
localparam signed [DEBIT:0]  W_6_x358 =  23'd32;
localparam signed [DEBIT:0]  W_6_x359 =  23'd189;
localparam signed [DEBIT:0]  W_6_x360 =  23'd453;
localparam signed [DEBIT:0]  W_6_x361 =  23'd656;
localparam signed [DEBIT:0]  W_6_x362 =  23'd806;
localparam signed [DEBIT:0]  W_6_x363 =  23'd906;
localparam signed [DEBIT:0]  W_6_x364 =  23'd967;
localparam signed [DEBIT:0]  W_6_x365 =  23'd963;
localparam signed [DEBIT:0]  W_6_x366 =  23'd964;
localparam signed [DEBIT:0]  W_6_x367 =  23'd929;
localparam signed [DEBIT:0]  W_6_x368 =  23'd801;
localparam signed [DEBIT:0]  W_6_x369 =  23'd517;
localparam signed [DEBIT:0]  W_6_x370 =  23'd125;
localparam signed [DEBIT:0]  W_6_x371 = - 23'd12;
localparam signed [DEBIT:0]  W_6_x372 =  23'd114;
localparam signed [DEBIT:0]  W_6_x373 =  23'd226;
localparam signed [DEBIT:0]  W_6_x374 =  23'd194;
localparam signed [DEBIT:0]  W_6_x375 =  23'd184;
localparam signed [DEBIT:0]  W_6_x376 =  23'd209;
localparam signed [DEBIT:0]  W_6_x377 =  23'd310;
localparam signed [DEBIT:0]  W_6_x378 = - 23'd80;
localparam signed [DEBIT:0]  W_6_x379 = - 23'd181;
localparam signed [DEBIT:0]  W_6_x380 =  23'd30;
localparam signed [DEBIT:0]  W_6_x381 =  23'd59;
localparam signed [DEBIT:0]  W_6_x382 = - 23'd50;
localparam signed [DEBIT:0]  W_6_x383 = - 23'd121;
localparam signed [DEBIT:0]  W_6_x384 = - 23'd105;
localparam signed [DEBIT:0]  W_6_x385 = - 23'd28;
localparam signed [DEBIT:0]  W_6_x386 =  23'd194;
localparam signed [DEBIT:0]  W_6_x387 =  23'd333;
localparam signed [DEBIT:0]  W_6_x388 =  23'd526;
localparam signed [DEBIT:0]  W_6_x389 =  23'd700;
localparam signed [DEBIT:0]  W_6_x390 =  23'd843;
localparam signed [DEBIT:0]  W_6_x391 =  23'd912;
localparam signed [DEBIT:0]  W_6_x392 =  23'd949;
localparam signed [DEBIT:0]  W_6_x393 =  23'd974;
localparam signed [DEBIT:0]  W_6_x394 =  23'd959;
localparam signed [DEBIT:0]  W_6_x395 =  23'd956;
localparam signed [DEBIT:0]  W_6_x396 =  23'd851;
localparam signed [DEBIT:0]  W_6_x397 =  23'd585;
localparam signed [DEBIT:0]  W_6_x398 =  23'd181;
localparam signed [DEBIT:0]  W_6_x399 =  23'd32;
localparam signed [DEBIT:0]  W_6_x400 =  23'd111;
localparam signed [DEBIT:0]  W_6_x401 =  23'd122;
localparam signed [DEBIT:0]  W_6_x402 =  23'd167;
localparam signed [DEBIT:0]  W_6_x403 =  23'd202;
localparam signed [DEBIT:0]  W_6_x404 =  23'd213;
localparam signed [DEBIT:0]  W_6_x405 =  23'd35;
localparam signed [DEBIT:0]  W_6_x406 = - 23'd305;
localparam signed [DEBIT:0]  W_6_x407 = - 23'd75;
localparam signed [DEBIT:0]  W_6_x408 =  23'd100;
localparam signed [DEBIT:0]  W_6_x409 =  23'd29;
localparam signed [DEBIT:0]  W_6_x410 = - 23'd147;
localparam signed [DEBIT:0]  W_6_x411 = - 23'd276;
localparam signed [DEBIT:0]  W_6_x412 = - 23'd157;
localparam signed [DEBIT:0]  W_6_x413 =  23'd30;
localparam signed [DEBIT:0]  W_6_x414 =  23'd294;
localparam signed [DEBIT:0]  W_6_x415 =  23'd391;
localparam signed [DEBIT:0]  W_6_x416 =  23'd447;
localparam signed [DEBIT:0]  W_6_x417 =  23'd666;
localparam signed [DEBIT:0]  W_6_x418 =  23'd878;
localparam signed [DEBIT:0]  W_6_x419 =  23'd918;
localparam signed [DEBIT:0]  W_6_x420 =  23'd974;
localparam signed [DEBIT:0]  W_6_x421 =  23'd969;
localparam signed [DEBIT:0]  W_6_x422 =  23'd965;
localparam signed [DEBIT:0]  W_6_x423 =  23'd966;
localparam signed [DEBIT:0]  W_6_x424 =  23'd860;
localparam signed [DEBIT:0]  W_6_x425 =  23'd584;
localparam signed [DEBIT:0]  W_6_x426 =  23'd124;
localparam signed [DEBIT:0]  W_6_x427 = - 23'd78;
localparam signed [DEBIT:0]  W_6_x428 =  23'd32;
localparam signed [DEBIT:0]  W_6_x429 =  23'd52;
localparam signed [DEBIT:0]  W_6_x430 =  23'd133;
localparam signed [DEBIT:0]  W_6_x431 =  23'd157;
localparam signed [DEBIT:0]  W_6_x432 =  23'd114;
localparam signed [DEBIT:0]  W_6_x433 = - 23'd13;
localparam signed [DEBIT:0]  W_6_x434 = - 23'd197;
localparam signed [DEBIT:0]  W_6_x435 =  23'd25;
localparam signed [DEBIT:0]  W_6_x436 =  23'd150;
localparam signed [DEBIT:0]  W_6_x437 = - 23'd3;
localparam signed [DEBIT:0]  W_6_x438 = - 23'd156;
localparam signed [DEBIT:0]  W_6_x439 = - 23'd214;
localparam signed [DEBIT:0]  W_6_x440 = - 23'd113;
localparam signed [DEBIT:0]  W_6_x441 =  23'd106;
localparam signed [DEBIT:0]  W_6_x442 =  23'd236;
localparam signed [DEBIT:0]  W_6_x443 =  23'd297;
localparam signed [DEBIT:0]  W_6_x444 =  23'd350;
localparam signed [DEBIT:0]  W_6_x445 =  23'd560;
localparam signed [DEBIT:0]  W_6_x446 =  23'd793;
localparam signed [DEBIT:0]  W_6_x447 =  23'd866;
localparam signed [DEBIT:0]  W_6_x448 =  23'd962;
localparam signed [DEBIT:0]  W_6_x449 =  23'd970;
localparam signed [DEBIT:0]  W_6_x450 =  23'd967;
localparam signed [DEBIT:0]  W_6_x451 =  23'd968;
localparam signed [DEBIT:0]  W_6_x452 =  23'd863;
localparam signed [DEBIT:0]  W_6_x453 =  23'd540;
localparam signed [DEBIT:0]  W_6_x454 = - 23'd15;
localparam signed [DEBIT:0]  W_6_x455 = - 23'd176;
localparam signed [DEBIT:0]  W_6_x456 =  23'd0;
localparam signed [DEBIT:0]  W_6_x457 =  23'd77;
localparam signed [DEBIT:0]  W_6_x458 =  23'd111;
localparam signed [DEBIT:0]  W_6_x459 =  23'd133;
localparam signed [DEBIT:0]  W_6_x460 =  23'd86;
localparam signed [DEBIT:0]  W_6_x461 = - 23'd63;
localparam signed [DEBIT:0]  W_6_x462 = - 23'd73;
localparam signed [DEBIT:0]  W_6_x463 =  23'd32;
localparam signed [DEBIT:0]  W_6_x464 = - 23'd73;
localparam signed [DEBIT:0]  W_6_x465 = - 23'd284;
localparam signed [DEBIT:0]  W_6_x466 = - 23'd235;
localparam signed [DEBIT:0]  W_6_x467 = - 23'd123;
localparam signed [DEBIT:0]  W_6_x468 =  23'd5;
localparam signed [DEBIT:0]  W_6_x469 =  23'd81;
localparam signed [DEBIT:0]  W_6_x470 =  23'd20;
localparam signed [DEBIT:0]  W_6_x471 =  23'd178;
localparam signed [DEBIT:0]  W_6_x472 =  23'd219;
localparam signed [DEBIT:0]  W_6_x473 =  23'd389;
localparam signed [DEBIT:0]  W_6_x474 =  23'd654;
localparam signed [DEBIT:0]  W_6_x475 =  23'd845;
localparam signed [DEBIT:0]  W_6_x476 =  23'd959;
localparam signed [DEBIT:0]  W_6_x477 =  23'd979;
localparam signed [DEBIT:0]  W_6_x478 =  23'd977;
localparam signed [DEBIT:0]  W_6_x479 =  23'd968;
localparam signed [DEBIT:0]  W_6_x480 =  23'd851;
localparam signed [DEBIT:0]  W_6_x481 =  23'd421;
localparam signed [DEBIT:0]  W_6_x482 = - 23'd132;
localparam signed [DEBIT:0]  W_6_x483 = - 23'd172;
localparam signed [DEBIT:0]  W_6_x484 =  23'd7;
localparam signed [DEBIT:0]  W_6_x485 =  23'd190;
localparam signed [DEBIT:0]  W_6_x486 =  23'd189;
localparam signed [DEBIT:0]  W_6_x487 =  23'd303;
localparam signed [DEBIT:0]  W_6_x488 =  23'd168;
localparam signed [DEBIT:0]  W_6_x489 =  23'd78;
localparam signed [DEBIT:0]  W_6_x490 = - 23'd48;
localparam signed [DEBIT:0]  W_6_x491 = - 23'd143;
localparam signed [DEBIT:0]  W_6_x492 = - 23'd322;
localparam signed [DEBIT:0]  W_6_x493 = - 23'd314;
localparam signed [DEBIT:0]  W_6_x494 = - 23'd125;
localparam signed [DEBIT:0]  W_6_x495 = - 23'd25;
localparam signed [DEBIT:0]  W_6_x496 =  23'd63;
localparam signed [DEBIT:0]  W_6_x497 =  23'd6;
localparam signed [DEBIT:0]  W_6_x498 = - 23'd102;
localparam signed [DEBIT:0]  W_6_x499 =  23'd21;
localparam signed [DEBIT:0]  W_6_x500 =  23'd82;
localparam signed [DEBIT:0]  W_6_x501 =  23'd251;
localparam signed [DEBIT:0]  W_6_x502 =  23'd593;
localparam signed [DEBIT:0]  W_6_x503 =  23'd846;
localparam signed [DEBIT:0]  W_6_x504 =  23'd961;
localparam signed [DEBIT:0]  W_6_x505 =  23'd969;
localparam signed [DEBIT:0]  W_6_x506 =  23'd974;
localparam signed [DEBIT:0]  W_6_x507 =  23'd970;
localparam signed [DEBIT:0]  W_6_x508 =  23'd807;
localparam signed [DEBIT:0]  W_6_x509 =  23'd327;
localparam signed [DEBIT:0]  W_6_x510 = - 23'd276;
localparam signed [DEBIT:0]  W_6_x511 = - 23'd286;
localparam signed [DEBIT:0]  W_6_x512 = - 23'd30;
localparam signed [DEBIT:0]  W_6_x513 =  23'd249;
localparam signed [DEBIT:0]  W_6_x514 =  23'd363;
localparam signed [DEBIT:0]  W_6_x515 =  23'd383;
localparam signed [DEBIT:0]  W_6_x516 =  23'd397;
localparam signed [DEBIT:0]  W_6_x517 =  23'd290;
localparam signed [DEBIT:0]  W_6_x518 = - 23'd5;
localparam signed [DEBIT:0]  W_6_x519 = - 23'd151;
localparam signed [DEBIT:0]  W_6_x520 = - 23'd151;
localparam signed [DEBIT:0]  W_6_x521 = - 23'd46;
localparam signed [DEBIT:0]  W_6_x522 = - 23'd46;
localparam signed [DEBIT:0]  W_6_x523 =  23'd85;
localparam signed [DEBIT:0]  W_6_x524 =  23'd34;
localparam signed [DEBIT:0]  W_6_x525 = - 23'd80;
localparam signed [DEBIT:0]  W_6_x526 = - 23'd127;
localparam signed [DEBIT:0]  W_6_x527 = - 23'd216;
localparam signed [DEBIT:0]  W_6_x528 = - 23'd71;
localparam signed [DEBIT:0]  W_6_x529 =  23'd223;
localparam signed [DEBIT:0]  W_6_x530 =  23'd669;
localparam signed [DEBIT:0]  W_6_x531 =  23'd885;
localparam signed [DEBIT:0]  W_6_x532 =  23'd972;
localparam signed [DEBIT:0]  W_6_x533 =  23'd967;
localparam signed [DEBIT:0]  W_6_x534 =  23'd961;
localparam signed [DEBIT:0]  W_6_x535 =  23'd951;
localparam signed [DEBIT:0]  W_6_x536 =  23'd747;
localparam signed [DEBIT:0]  W_6_x537 =  23'd247;
localparam signed [DEBIT:0]  W_6_x538 = - 23'd279;
localparam signed [DEBIT:0]  W_6_x539 = - 23'd495;
localparam signed [DEBIT:0]  W_6_x540 = - 23'd284;
localparam signed [DEBIT:0]  W_6_x541 = - 23'd32;
localparam signed [DEBIT:0]  W_6_x542 =  23'd194;
localparam signed [DEBIT:0]  W_6_x543 =  23'd366;
localparam signed [DEBIT:0]  W_6_x544 =  23'd441;
localparam signed [DEBIT:0]  W_6_x545 =  23'd338;
localparam signed [DEBIT:0]  W_6_x546 =  23'd106;
localparam signed [DEBIT:0]  W_6_x547 =  23'd63;
localparam signed [DEBIT:0]  W_6_x548 =  23'd151;
localparam signed [DEBIT:0]  W_6_x549 =  23'd137;
localparam signed [DEBIT:0]  W_6_x550 =  23'd42;
localparam signed [DEBIT:0]  W_6_x551 = - 23'd52;
localparam signed [DEBIT:0]  W_6_x552 = - 23'd158;
localparam signed [DEBIT:0]  W_6_x553 = - 23'd206;
localparam signed [DEBIT:0]  W_6_x554 = - 23'd358;
localparam signed [DEBIT:0]  W_6_x555 = - 23'd416;
localparam signed [DEBIT:0]  W_6_x556 = - 23'd138;
localparam signed [DEBIT:0]  W_6_x557 =  23'd349;
localparam signed [DEBIT:0]  W_6_x558 =  23'd744;
localparam signed [DEBIT:0]  W_6_x559 =  23'd920;
localparam signed [DEBIT:0]  W_6_x560 =  23'd968;
localparam signed [DEBIT:0]  W_6_x561 =  23'd972;
localparam signed [DEBIT:0]  W_6_x562 =  23'd968;
localparam signed [DEBIT:0]  W_6_x563 =  23'd940;
localparam signed [DEBIT:0]  W_6_x564 =  23'd710;
localparam signed [DEBIT:0]  W_6_x565 =  23'd224;
localparam signed [DEBIT:0]  W_6_x566 = - 23'd247;
localparam signed [DEBIT:0]  W_6_x567 = - 23'd530;
localparam signed [DEBIT:0]  W_6_x568 = - 23'd400;
localparam signed [DEBIT:0]  W_6_x569 = - 23'd306;
localparam signed [DEBIT:0]  W_6_x570 = - 23'd126;
localparam signed [DEBIT:0]  W_6_x571 =  23'd157;
localparam signed [DEBIT:0]  W_6_x572 =  23'd229;
localparam signed [DEBIT:0]  W_6_x573 =  23'd261;
localparam signed [DEBIT:0]  W_6_x574 =  23'd254;
localparam signed [DEBIT:0]  W_6_x575 =  23'd283;
localparam signed [DEBIT:0]  W_6_x576 =  23'd209;
localparam signed [DEBIT:0]  W_6_x577 =  23'd125;
localparam signed [DEBIT:0]  W_6_x578 =  23'd39;
localparam signed [DEBIT:0]  W_6_x579 = - 23'd72;
localparam signed [DEBIT:0]  W_6_x580 = - 23'd278;
localparam signed [DEBIT:0]  W_6_x581 = - 23'd414;
localparam signed [DEBIT:0]  W_6_x582 = - 23'd460;
localparam signed [DEBIT:0]  W_6_x583 = - 23'd452;
localparam signed [DEBIT:0]  W_6_x584 = - 23'd9;
localparam signed [DEBIT:0]  W_6_x585 =  23'd510;
localparam signed [DEBIT:0]  W_6_x586 =  23'd823;
localparam signed [DEBIT:0]  W_6_x587 =  23'd960;
localparam signed [DEBIT:0]  W_6_x588 =  23'd972;
localparam signed [DEBIT:0]  W_6_x589 =  23'd972;
localparam signed [DEBIT:0]  W_6_x590 =  23'd972;
localparam signed [DEBIT:0]  W_6_x591 =  23'd947;
localparam signed [DEBIT:0]  W_6_x592 =  23'd792;
localparam signed [DEBIT:0]  W_6_x593 =  23'd354;
localparam signed [DEBIT:0]  W_6_x594 = - 23'd84;
localparam signed [DEBIT:0]  W_6_x595 = - 23'd443;
localparam signed [DEBIT:0]  W_6_x596 = - 23'd540;
localparam signed [DEBIT:0]  W_6_x597 = - 23'd428;
localparam signed [DEBIT:0]  W_6_x598 = - 23'd333;
localparam signed [DEBIT:0]  W_6_x599 = - 23'd29;
localparam signed [DEBIT:0]  W_6_x600 =  23'd197;
localparam signed [DEBIT:0]  W_6_x601 =  23'd328;
localparam signed [DEBIT:0]  W_6_x602 =  23'd428;
localparam signed [DEBIT:0]  W_6_x603 =  23'd411;
localparam signed [DEBIT:0]  W_6_x604 =  23'd286;
localparam signed [DEBIT:0]  W_6_x605 =  23'd192;
localparam signed [DEBIT:0]  W_6_x606 =  23'd176;
localparam signed [DEBIT:0]  W_6_x607 =  23'd19;
localparam signed [DEBIT:0]  W_6_x608 = - 23'd282;
localparam signed [DEBIT:0]  W_6_x609 = - 23'd496;
localparam signed [DEBIT:0]  W_6_x610 = - 23'd448;
localparam signed [DEBIT:0]  W_6_x611 = - 23'd206;
localparam signed [DEBIT:0]  W_6_x612 =  23'd287;
localparam signed [DEBIT:0]  W_6_x613 =  23'd660;
localparam signed [DEBIT:0]  W_6_x614 =  23'd894;
localparam signed [DEBIT:0]  W_6_x615 =  23'd958;
localparam signed [DEBIT:0]  W_6_x616 =  23'd977;
localparam signed [DEBIT:0]  W_6_x617 =  23'd969;
localparam signed [DEBIT:0]  W_6_x618 =  23'd969;
localparam signed [DEBIT:0]  W_6_x619 =  23'd958;
localparam signed [DEBIT:0]  W_6_x620 =  23'd876;
localparam signed [DEBIT:0]  W_6_x621 =  23'd638;
localparam signed [DEBIT:0]  W_6_x622 =  23'd274;
localparam signed [DEBIT:0]  W_6_x623 = - 23'd35;
localparam signed [DEBIT:0]  W_6_x624 = - 23'd281;
localparam signed [DEBIT:0]  W_6_x625 = - 23'd298;
localparam signed [DEBIT:0]  W_6_x626 = - 23'd286;
localparam signed [DEBIT:0]  W_6_x627 = - 23'd120;
localparam signed [DEBIT:0]  W_6_x628 = - 23'd78;
localparam signed [DEBIT:0]  W_6_x629 =  23'd57;
localparam signed [DEBIT:0]  W_6_x630 =  23'd83;
localparam signed [DEBIT:0]  W_6_x631 =  23'd95;
localparam signed [DEBIT:0]  W_6_x632 =  23'd153;
localparam signed [DEBIT:0]  W_6_x633 =  23'd85;
localparam signed [DEBIT:0]  W_6_x634 = - 23'd26;
localparam signed [DEBIT:0]  W_6_x635 = - 23'd189;
localparam signed [DEBIT:0]  W_6_x636 = - 23'd303;
localparam signed [DEBIT:0]  W_6_x637 = - 23'd285;
localparam signed [DEBIT:0]  W_6_x638 = - 23'd111;
localparam signed [DEBIT:0]  W_6_x639 =  23'd185;
localparam signed [DEBIT:0]  W_6_x640 =  23'd574;
localparam signed [DEBIT:0]  W_6_x641 =  23'd837;
localparam signed [DEBIT:0]  W_6_x642 =  23'd939;
localparam signed [DEBIT:0]  W_6_x643 =  23'd965;
localparam signed [DEBIT:0]  W_6_x644 =  23'd971;
localparam signed [DEBIT:0]  W_6_x645 =  23'd978;
localparam signed [DEBIT:0]  W_6_x646 =  23'd973;
localparam signed [DEBIT:0]  W_6_x647 =  23'd970;
localparam signed [DEBIT:0]  W_6_x648 =  23'd931;
localparam signed [DEBIT:0]  W_6_x649 =  23'd867;
localparam signed [DEBIT:0]  W_6_x650 =  23'd719;
localparam signed [DEBIT:0]  W_6_x651 =  23'd489;
localparam signed [DEBIT:0]  W_6_x652 =  23'd213;
localparam signed [DEBIT:0]  W_6_x653 =  23'd39;
localparam signed [DEBIT:0]  W_6_x654 = - 23'd105;
localparam signed [DEBIT:0]  W_6_x655 = - 23'd204;
localparam signed [DEBIT:0]  W_6_x656 = - 23'd191;
localparam signed [DEBIT:0]  W_6_x657 = - 23'd150;
localparam signed [DEBIT:0]  W_6_x658 = - 23'd122;
localparam signed [DEBIT:0]  W_6_x659 = - 23'd137;
localparam signed [DEBIT:0]  W_6_x660 = - 23'd52;
localparam signed [DEBIT:0]  W_6_x661 = - 23'd49;
localparam signed [DEBIT:0]  W_6_x662 = - 23'd70;
localparam signed [DEBIT:0]  W_6_x663 = - 23'd23;
localparam signed [DEBIT:0]  W_6_x664 =  23'd94;
localparam signed [DEBIT:0]  W_6_x665 =  23'd187;
localparam signed [DEBIT:0]  W_6_x666 =  23'd366;
localparam signed [DEBIT:0]  W_6_x667 =  23'd584;
localparam signed [DEBIT:0]  W_6_x668 =  23'd786;
localparam signed [DEBIT:0]  W_6_x669 =  23'd923;
localparam signed [DEBIT:0]  W_6_x670 =  23'd973;
localparam signed [DEBIT:0]  W_6_x671 =  23'd970;
localparam signed [DEBIT:0]  W_6_x672 =  23'd969;
localparam signed [DEBIT:0]  W_6_x673 =  23'd976;
localparam signed [DEBIT:0]  W_6_x674 =  23'd965;
localparam signed [DEBIT:0]  W_6_x675 =  23'd981;
localparam signed [DEBIT:0]  W_6_x676 =  23'd959;
localparam signed [DEBIT:0]  W_6_x677 =  23'd926;
localparam signed [DEBIT:0]  W_6_x678 =  23'd881;
localparam signed [DEBIT:0]  W_6_x679 =  23'd801;
localparam signed [DEBIT:0]  W_6_x680 =  23'd647;
localparam signed [DEBIT:0]  W_6_x681 =  23'd504;
localparam signed [DEBIT:0]  W_6_x682 =  23'd319;
localparam signed [DEBIT:0]  W_6_x683 =  23'd217;
localparam signed [DEBIT:0]  W_6_x684 =  23'd242;
localparam signed [DEBIT:0]  W_6_x685 =  23'd292;
localparam signed [DEBIT:0]  W_6_x686 =  23'd199;
localparam signed [DEBIT:0]  W_6_x687 =  23'd157;
localparam signed [DEBIT:0]  W_6_x688 =  23'd153;
localparam signed [DEBIT:0]  W_6_x689 =  23'd153;
localparam signed [DEBIT:0]  W_6_x690 =  23'd196;
localparam signed [DEBIT:0]  W_6_x691 =  23'd290;
localparam signed [DEBIT:0]  W_6_x692 =  23'd438;
localparam signed [DEBIT:0]  W_6_x693 =  23'd521;
localparam signed [DEBIT:0]  W_6_x694 =  23'd646;
localparam signed [DEBIT:0]  W_6_x695 =  23'd765;
localparam signed [DEBIT:0]  W_6_x696 =  23'd887;
localparam signed [DEBIT:0]  W_6_x697 =  23'd955;
localparam signed [DEBIT:0]  W_6_x698 =  23'd965;
localparam signed [DEBIT:0]  W_6_x699 =  23'd973;
localparam signed [DEBIT:0]  W_6_x700 =  23'd974;
localparam signed [DEBIT:0]  W_6_x701 =  23'd974;
localparam signed [DEBIT:0]  W_6_x702 =  23'd968;
localparam signed [DEBIT:0]  W_6_x703 =  23'd970;
localparam signed [DEBIT:0]  W_6_x704 =  23'd971;
localparam signed [DEBIT:0]  W_6_x705 =  23'd958;
localparam signed [DEBIT:0]  W_6_x706 =  23'd959;
localparam signed [DEBIT:0]  W_6_x707 =  23'd923;
localparam signed [DEBIT:0]  W_6_x708 =  23'd873;
localparam signed [DEBIT:0]  W_6_x709 =  23'd806;
localparam signed [DEBIT:0]  W_6_x710 =  23'd708;
localparam signed [DEBIT:0]  W_6_x711 =  23'd671;
localparam signed [DEBIT:0]  W_6_x712 =  23'd698;
localparam signed [DEBIT:0]  W_6_x713 =  23'd645;
localparam signed [DEBIT:0]  W_6_x714 =  23'd594;
localparam signed [DEBIT:0]  W_6_x715 =  23'd552;
localparam signed [DEBIT:0]  W_6_x716 =  23'd567;
localparam signed [DEBIT:0]  W_6_x717 =  23'd526;
localparam signed [DEBIT:0]  W_6_x718 =  23'd569;
localparam signed [DEBIT:0]  W_6_x719 =  23'd625;
localparam signed [DEBIT:0]  W_6_x720 =  23'd704;
localparam signed [DEBIT:0]  W_6_x721 =  23'd757;
localparam signed [DEBIT:0]  W_6_x722 =  23'd829;
localparam signed [DEBIT:0]  W_6_x723 =  23'd881;
localparam signed [DEBIT:0]  W_6_x724 =  23'd936;
localparam signed [DEBIT:0]  W_6_x725 =  23'd959;
localparam signed [DEBIT:0]  W_6_x726 =  23'd967;
localparam signed [DEBIT:0]  W_6_x727 =  23'd975;
localparam signed [DEBIT:0]  W_6_x728 =  23'd976;
localparam signed [DEBIT:0]  W_6_x729 =  23'd976;
localparam signed [DEBIT:0]  W_6_x730 =  23'd974;
localparam signed [DEBIT:0]  W_6_x731 =  23'd954;
localparam signed [DEBIT:0]  W_6_x732 =  23'd972;
localparam signed [DEBIT:0]  W_6_x733 =  23'd965;
localparam signed [DEBIT:0]  W_6_x734 =  23'd948;
localparam signed [DEBIT:0]  W_6_x735 =  23'd935;
localparam signed [DEBIT:0]  W_6_x736 =  23'd927;
localparam signed [DEBIT:0]  W_6_x737 =  23'd900;
localparam signed [DEBIT:0]  W_6_x738 =  23'd881;
localparam signed [DEBIT:0]  W_6_x739 =  23'd869;
localparam signed [DEBIT:0]  W_6_x740 =  23'd877;
localparam signed [DEBIT:0]  W_6_x741 =  23'd868;
localparam signed [DEBIT:0]  W_6_x742 =  23'd829;
localparam signed [DEBIT:0]  W_6_x743 =  23'd787;
localparam signed [DEBIT:0]  W_6_x744 =  23'd774;
localparam signed [DEBIT:0]  W_6_x745 =  23'd738;
localparam signed [DEBIT:0]  W_6_x746 =  23'd737;
localparam signed [DEBIT:0]  W_6_x747 =  23'd772;
localparam signed [DEBIT:0]  W_6_x748 =  23'd832;
localparam signed [DEBIT:0]  W_6_x749 =  23'd882;
localparam signed [DEBIT:0]  W_6_x750 =  23'd890;
localparam signed [DEBIT:0]  W_6_x751 =  23'd930;
localparam signed [DEBIT:0]  W_6_x752 =  23'd966;
localparam signed [DEBIT:0]  W_6_x753 =  23'd970;
localparam signed [DEBIT:0]  W_6_x754 =  23'd968;
localparam signed [DEBIT:0]  W_6_x755 =  23'd967;
localparam signed [DEBIT:0]  W_6_x756 =  23'd973;
localparam signed [DEBIT:0]  W_6_x757 =  23'd967;
localparam signed [DEBIT:0]  W_6_x758 =  23'd970;
localparam signed [DEBIT:0]  W_6_x759 =  23'd964;
localparam signed [DEBIT:0]  W_6_x760 =  23'd968;
localparam signed [DEBIT:0]  W_6_x761 =  23'd975;
localparam signed [DEBIT:0]  W_6_x762 =  23'd957;
localparam signed [DEBIT:0]  W_6_x763 =  23'd953;
localparam signed [DEBIT:0]  W_6_x764 =  23'd927;
localparam signed [DEBIT:0]  W_6_x765 =  23'd965;
localparam signed [DEBIT:0]  W_6_x766 =  23'd978;
localparam signed [DEBIT:0]  W_6_x767 =  23'd971;
localparam signed [DEBIT:0]  W_6_x768 =  23'd954;
localparam signed [DEBIT:0]  W_6_x769 =  23'd935;
localparam signed [DEBIT:0]  W_6_x770 =  23'd941;
localparam signed [DEBIT:0]  W_6_x771 =  23'd919;
localparam signed [DEBIT:0]  W_6_x772 =  23'd915;
localparam signed [DEBIT:0]  W_6_x773 =  23'd895;
localparam signed [DEBIT:0]  W_6_x774 =  23'd884;
localparam signed [DEBIT:0]  W_6_x775 =  23'd892;
localparam signed [DEBIT:0]  W_6_x776 =  23'd927;
localparam signed [DEBIT:0]  W_6_x777 =  23'd953;
localparam signed [DEBIT:0]  W_6_x778 =  23'd954;
localparam signed [DEBIT:0]  W_6_x779 =  23'd969;
localparam signed [DEBIT:0]  W_6_x780 =  23'd967;
localparam signed [DEBIT:0]  W_6_x781 =  23'd965;
localparam signed [DEBIT:0]  W_6_x782 =  23'd974;
localparam signed [DEBIT:0]  W_6_x783 =  23'd972;
localparam signed [DEBIT:0]  W_6_x784 =  23'd974;
localparam signed [DEBIT:0]  W_7_x1 =  23'd972;
localparam signed [DEBIT:0]  W_7_x2 =  23'd988;
localparam signed [DEBIT:0]  W_7_x3 =  23'd976;
localparam signed [DEBIT:0]  W_7_x4 =  23'd975;
localparam signed [DEBIT:0]  W_7_x5 =  23'd970;
localparam signed [DEBIT:0]  W_7_x6 =  23'd980;
localparam signed [DEBIT:0]  W_7_x7 =  23'd981;
localparam signed [DEBIT:0]  W_7_x8 =  23'd972;
localparam signed [DEBIT:0]  W_7_x9 =  23'd990;
localparam signed [DEBIT:0]  W_7_x10 =  23'd982;
localparam signed [DEBIT:0]  W_7_x11 =  23'd976;
localparam signed [DEBIT:0]  W_7_x12 =  23'd985;
localparam signed [DEBIT:0]  W_7_x13 =  23'd979;
localparam signed [DEBIT:0]  W_7_x14 =  23'd977;
localparam signed [DEBIT:0]  W_7_x15 =  23'd976;
localparam signed [DEBIT:0]  W_7_x16 =  23'd969;
localparam signed [DEBIT:0]  W_7_x17 =  23'd979;
localparam signed [DEBIT:0]  W_7_x18 =  23'd981;
localparam signed [DEBIT:0]  W_7_x19 =  23'd972;
localparam signed [DEBIT:0]  W_7_x20 =  23'd975;
localparam signed [DEBIT:0]  W_7_x21 =  23'd979;
localparam signed [DEBIT:0]  W_7_x22 =  23'd976;
localparam signed [DEBIT:0]  W_7_x23 =  23'd977;
localparam signed [DEBIT:0]  W_7_x24 =  23'd977;
localparam signed [DEBIT:0]  W_7_x25 =  23'd990;
localparam signed [DEBIT:0]  W_7_x26 =  23'd984;
localparam signed [DEBIT:0]  W_7_x27 =  23'd972;
localparam signed [DEBIT:0]  W_7_x28 =  23'd976;
localparam signed [DEBIT:0]  W_7_x29 =  23'd978;
localparam signed [DEBIT:0]  W_7_x30 =  23'd988;
localparam signed [DEBIT:0]  W_7_x31 =  23'd970;
localparam signed [DEBIT:0]  W_7_x32 =  23'd977;
localparam signed [DEBIT:0]  W_7_x33 =  23'd972;
localparam signed [DEBIT:0]  W_7_x34 =  23'd975;
localparam signed [DEBIT:0]  W_7_x35 =  23'd976;
localparam signed [DEBIT:0]  W_7_x36 =  23'd978;
localparam signed [DEBIT:0]  W_7_x37 =  23'd965;
localparam signed [DEBIT:0]  W_7_x38 =  23'd952;
localparam signed [DEBIT:0]  W_7_x39 =  23'd962;
localparam signed [DEBIT:0]  W_7_x40 =  23'd970;
localparam signed [DEBIT:0]  W_7_x41 =  23'd947;
localparam signed [DEBIT:0]  W_7_x42 =  23'd950;
localparam signed [DEBIT:0]  W_7_x43 =  23'd942;
localparam signed [DEBIT:0]  W_7_x44 =  23'd953;
localparam signed [DEBIT:0]  W_7_x45 =  23'd959;
localparam signed [DEBIT:0]  W_7_x46 =  23'd976;
localparam signed [DEBIT:0]  W_7_x47 =  23'd969;
localparam signed [DEBIT:0]  W_7_x48 =  23'd965;
localparam signed [DEBIT:0]  W_7_x49 =  23'd974;
localparam signed [DEBIT:0]  W_7_x50 =  23'd981;
localparam signed [DEBIT:0]  W_7_x51 =  23'd982;
localparam signed [DEBIT:0]  W_7_x52 =  23'd969;
localparam signed [DEBIT:0]  W_7_x53 =  23'd976;
localparam signed [DEBIT:0]  W_7_x54 =  23'd982;
localparam signed [DEBIT:0]  W_7_x55 =  23'd979;
localparam signed [DEBIT:0]  W_7_x56 =  23'd988;
localparam signed [DEBIT:0]  W_7_x57 =  23'd980;
localparam signed [DEBIT:0]  W_7_x58 =  23'd986;
localparam signed [DEBIT:0]  W_7_x59 =  23'd976;
localparam signed [DEBIT:0]  W_7_x60 =  23'd979;
localparam signed [DEBIT:0]  W_7_x61 =  23'd980;
localparam signed [DEBIT:0]  W_7_x62 =  23'd983;
localparam signed [DEBIT:0]  W_7_x63 =  23'd963;
localparam signed [DEBIT:0]  W_7_x64 =  23'd939;
localparam signed [DEBIT:0]  W_7_x65 =  23'd908;
localparam signed [DEBIT:0]  W_7_x66 =  23'd875;
localparam signed [DEBIT:0]  W_7_x67 =  23'd866;
localparam signed [DEBIT:0]  W_7_x68 =  23'd875;
localparam signed [DEBIT:0]  W_7_x69 =  23'd841;
localparam signed [DEBIT:0]  W_7_x70 =  23'd831;
localparam signed [DEBIT:0]  W_7_x71 =  23'd803;
localparam signed [DEBIT:0]  W_7_x72 =  23'd819;
localparam signed [DEBIT:0]  W_7_x73 =  23'd837;
localparam signed [DEBIT:0]  W_7_x74 =  23'd889;
localparam signed [DEBIT:0]  W_7_x75 =  23'd922;
localparam signed [DEBIT:0]  W_7_x76 =  23'd954;
localparam signed [DEBIT:0]  W_7_x77 =  23'd978;
localparam signed [DEBIT:0]  W_7_x78 =  23'd978;
localparam signed [DEBIT:0]  W_7_x79 =  23'd977;
localparam signed [DEBIT:0]  W_7_x80 =  23'd970;
localparam signed [DEBIT:0]  W_7_x81 =  23'd986;
localparam signed [DEBIT:0]  W_7_x82 =  23'd983;
localparam signed [DEBIT:0]  W_7_x83 =  23'd992;
localparam signed [DEBIT:0]  W_7_x84 =  23'd976;
localparam signed [DEBIT:0]  W_7_x85 =  23'd976;
localparam signed [DEBIT:0]  W_7_x86 =  23'd980;
localparam signed [DEBIT:0]  W_7_x87 =  23'd975;
localparam signed [DEBIT:0]  W_7_x88 =  23'd975;
localparam signed [DEBIT:0]  W_7_x89 =  23'd971;
localparam signed [DEBIT:0]  W_7_x90 =  23'd965;
localparam signed [DEBIT:0]  W_7_x91 =  23'd927;
localparam signed [DEBIT:0]  W_7_x92 =  23'd850;
localparam signed [DEBIT:0]  W_7_x93 =  23'd750;
localparam signed [DEBIT:0]  W_7_x94 =  23'd700;
localparam signed [DEBIT:0]  W_7_x95 =  23'd626;
localparam signed [DEBIT:0]  W_7_x96 =  23'd556;
localparam signed [DEBIT:0]  W_7_x97 =  23'd508;
localparam signed [DEBIT:0]  W_7_x98 =  23'd524;
localparam signed [DEBIT:0]  W_7_x99 =  23'd528;
localparam signed [DEBIT:0]  W_7_x100 =  23'd517;
localparam signed [DEBIT:0]  W_7_x101 =  23'd540;
localparam signed [DEBIT:0]  W_7_x102 =  23'd625;
localparam signed [DEBIT:0]  W_7_x103 =  23'd690;
localparam signed [DEBIT:0]  W_7_x104 =  23'd774;
localparam signed [DEBIT:0]  W_7_x105 =  23'd838;
localparam signed [DEBIT:0]  W_7_x106 =  23'd899;
localparam signed [DEBIT:0]  W_7_x107 =  23'd947;
localparam signed [DEBIT:0]  W_7_x108 =  23'd963;
localparam signed [DEBIT:0]  W_7_x109 =  23'd975;
localparam signed [DEBIT:0]  W_7_x110 =  23'd977;
localparam signed [DEBIT:0]  W_7_x111 =  23'd981;
localparam signed [DEBIT:0]  W_7_x112 =  23'd975;
localparam signed [DEBIT:0]  W_7_x113 =  23'd978;
localparam signed [DEBIT:0]  W_7_x114 =  23'd976;
localparam signed [DEBIT:0]  W_7_x115 =  23'd978;
localparam signed [DEBIT:0]  W_7_x116 =  23'd985;
localparam signed [DEBIT:0]  W_7_x117 =  23'd967;
localparam signed [DEBIT:0]  W_7_x118 =  23'd909;
localparam signed [DEBIT:0]  W_7_x119 =  23'd807;
localparam signed [DEBIT:0]  W_7_x120 =  23'd676;
localparam signed [DEBIT:0]  W_7_x121 =  23'd507;
localparam signed [DEBIT:0]  W_7_x122 =  23'd376;
localparam signed [DEBIT:0]  W_7_x123 =  23'd331;
localparam signed [DEBIT:0]  W_7_x124 =  23'd289;
localparam signed [DEBIT:0]  W_7_x125 =  23'd181;
localparam signed [DEBIT:0]  W_7_x126 =  23'd166;
localparam signed [DEBIT:0]  W_7_x127 =  23'd163;
localparam signed [DEBIT:0]  W_7_x128 =  23'd59;
localparam signed [DEBIT:0]  W_7_x129 =  23'd35;
localparam signed [DEBIT:0]  W_7_x130 =  23'd133;
localparam signed [DEBIT:0]  W_7_x131 =  23'd252;
localparam signed [DEBIT:0]  W_7_x132 =  23'd363;
localparam signed [DEBIT:0]  W_7_x133 =  23'd483;
localparam signed [DEBIT:0]  W_7_x134 =  23'd670;
localparam signed [DEBIT:0]  W_7_x135 =  23'd775;
localparam signed [DEBIT:0]  W_7_x136 =  23'd889;
localparam signed [DEBIT:0]  W_7_x137 =  23'd956;
localparam signed [DEBIT:0]  W_7_x138 =  23'd979;
localparam signed [DEBIT:0]  W_7_x139 =  23'd983;
localparam signed [DEBIT:0]  W_7_x140 =  23'd1005;
localparam signed [DEBIT:0]  W_7_x141 =  23'd986;
localparam signed [DEBIT:0]  W_7_x142 =  23'd975;
localparam signed [DEBIT:0]  W_7_x143 =  23'd978;
localparam signed [DEBIT:0]  W_7_x144 =  23'd967;
localparam signed [DEBIT:0]  W_7_x145 =  23'd925;
localparam signed [DEBIT:0]  W_7_x146 =  23'd759;
localparam signed [DEBIT:0]  W_7_x147 =  23'd496;
localparam signed [DEBIT:0]  W_7_x148 =  23'd311;
localparam signed [DEBIT:0]  W_7_x149 =  23'd139;
localparam signed [DEBIT:0]  W_7_x150 =  23'd92;
localparam signed [DEBIT:0]  W_7_x151 =  23'd14;
localparam signed [DEBIT:0]  W_7_x152 = - 23'd58;
localparam signed [DEBIT:0]  W_7_x153 = - 23'd95;
localparam signed [DEBIT:0]  W_7_x154 = - 23'd229;
localparam signed [DEBIT:0]  W_7_x155 = - 23'd215;
localparam signed [DEBIT:0]  W_7_x156 = - 23'd253;
localparam signed [DEBIT:0]  W_7_x157 = - 23'd271;
localparam signed [DEBIT:0]  W_7_x158 = - 23'd265;
localparam signed [DEBIT:0]  W_7_x159 = - 23'd213;
localparam signed [DEBIT:0]  W_7_x160 = - 23'd104;
localparam signed [DEBIT:0]  W_7_x161 =  23'd54;
localparam signed [DEBIT:0]  W_7_x162 =  23'd286;
localparam signed [DEBIT:0]  W_7_x163 =  23'd515;
localparam signed [DEBIT:0]  W_7_x164 =  23'd684;
localparam signed [DEBIT:0]  W_7_x165 =  23'd824;
localparam signed [DEBIT:0]  W_7_x166 =  23'd932;
localparam signed [DEBIT:0]  W_7_x167 =  23'd968;
localparam signed [DEBIT:0]  W_7_x168 =  23'd972;
localparam signed [DEBIT:0]  W_7_x169 =  23'd971;
localparam signed [DEBIT:0]  W_7_x170 =  23'd978;
localparam signed [DEBIT:0]  W_7_x171 =  23'd966;
localparam signed [DEBIT:0]  W_7_x172 =  23'd914;
localparam signed [DEBIT:0]  W_7_x173 =  23'd776;
localparam signed [DEBIT:0]  W_7_x174 =  23'd545;
localparam signed [DEBIT:0]  W_7_x175 =  23'd293;
localparam signed [DEBIT:0]  W_7_x176 =  23'd99;
localparam signed [DEBIT:0]  W_7_x177 =  23'd8;
localparam signed [DEBIT:0]  W_7_x178 = - 23'd61;
localparam signed [DEBIT:0]  W_7_x179 = - 23'd59;
localparam signed [DEBIT:0]  W_7_x180 =  23'd34;
localparam signed [DEBIT:0]  W_7_x181 = - 23'd5;
localparam signed [DEBIT:0]  W_7_x182 = - 23'd110;
localparam signed [DEBIT:0]  W_7_x183 = - 23'd112;
localparam signed [DEBIT:0]  W_7_x184 = - 23'd87;
localparam signed [DEBIT:0]  W_7_x185 =  23'd24;
localparam signed [DEBIT:0]  W_7_x186 =  23'd70;
localparam signed [DEBIT:0]  W_7_x187 = - 23'd91;
localparam signed [DEBIT:0]  W_7_x188 = - 23'd176;
localparam signed [DEBIT:0]  W_7_x189 = - 23'd239;
localparam signed [DEBIT:0]  W_7_x190 = - 23'd138;
localparam signed [DEBIT:0]  W_7_x191 =  23'd71;
localparam signed [DEBIT:0]  W_7_x192 =  23'd371;
localparam signed [DEBIT:0]  W_7_x193 =  23'd581;
localparam signed [DEBIT:0]  W_7_x194 =  23'd730;
localparam signed [DEBIT:0]  W_7_x195 =  23'd895;
localparam signed [DEBIT:0]  W_7_x196 =  23'd966;
localparam signed [DEBIT:0]  W_7_x197 =  23'd979;
localparam signed [DEBIT:0]  W_7_x198 =  23'd987;
localparam signed [DEBIT:0]  W_7_x199 =  23'd973;
localparam signed [DEBIT:0]  W_7_x200 =  23'd855;
localparam signed [DEBIT:0]  W_7_x201 =  23'd652;
localparam signed [DEBIT:0]  W_7_x202 =  23'd366;
localparam signed [DEBIT:0]  W_7_x203 =  23'd150;
localparam signed [DEBIT:0]  W_7_x204 =  23'd38;
localparam signed [DEBIT:0]  W_7_x205 =  23'd38;
localparam signed [DEBIT:0]  W_7_x206 =  23'd76;
localparam signed [DEBIT:0]  W_7_x207 =  23'd233;
localparam signed [DEBIT:0]  W_7_x208 =  23'd256;
localparam signed [DEBIT:0]  W_7_x209 =  23'd99;
localparam signed [DEBIT:0]  W_7_x210 = - 23'd167;
localparam signed [DEBIT:0]  W_7_x211 = - 23'd280;
localparam signed [DEBIT:0]  W_7_x212 = - 23'd270;
localparam signed [DEBIT:0]  W_7_x213 = - 23'd201;
localparam signed [DEBIT:0]  W_7_x214 = - 23'd26;
localparam signed [DEBIT:0]  W_7_x215 = - 23'd7;
localparam signed [DEBIT:0]  W_7_x216 = - 23'd44;
localparam signed [DEBIT:0]  W_7_x217 = - 23'd214;
localparam signed [DEBIT:0]  W_7_x218 = - 23'd292;
localparam signed [DEBIT:0]  W_7_x219 = - 23'd216;
localparam signed [DEBIT:0]  W_7_x220 =  23'd52;
localparam signed [DEBIT:0]  W_7_x221 =  23'd431;
localparam signed [DEBIT:0]  W_7_x222 =  23'd681;
localparam signed [DEBIT:0]  W_7_x223 =  23'd881;
localparam signed [DEBIT:0]  W_7_x224 =  23'd967;
localparam signed [DEBIT:0]  W_7_x225 =  23'd984;
localparam signed [DEBIT:0]  W_7_x226 =  23'd970;
localparam signed [DEBIT:0]  W_7_x227 =  23'd967;
localparam signed [DEBIT:0]  W_7_x228 =  23'd819;
localparam signed [DEBIT:0]  W_7_x229 =  23'd574;
localparam signed [DEBIT:0]  W_7_x230 =  23'd315;
localparam signed [DEBIT:0]  W_7_x231 =  23'd104;
localparam signed [DEBIT:0]  W_7_x232 =  23'd115;
localparam signed [DEBIT:0]  W_7_x233 =  23'd121;
localparam signed [DEBIT:0]  W_7_x234 =  23'd206;
localparam signed [DEBIT:0]  W_7_x235 =  23'd217;
localparam signed [DEBIT:0]  W_7_x236 =  23'd225;
localparam signed [DEBIT:0]  W_7_x237 =  23'd66;
localparam signed [DEBIT:0]  W_7_x238 = - 23'd106;
localparam signed [DEBIT:0]  W_7_x239 = - 23'd170;
localparam signed [DEBIT:0]  W_7_x240 = - 23'd77;
localparam signed [DEBIT:0]  W_7_x241 = - 23'd82;
localparam signed [DEBIT:0]  W_7_x242 = - 23'd45;
localparam signed [DEBIT:0]  W_7_x243 = - 23'd75;
localparam signed [DEBIT:0]  W_7_x244 = - 23'd1;
localparam signed [DEBIT:0]  W_7_x245 = - 23'd114;
localparam signed [DEBIT:0]  W_7_x246 = - 23'd325;
localparam signed [DEBIT:0]  W_7_x247 = - 23'd172;
localparam signed [DEBIT:0]  W_7_x248 =  23'd43;
localparam signed [DEBIT:0]  W_7_x249 =  23'd443;
localparam signed [DEBIT:0]  W_7_x250 =  23'd697;
localparam signed [DEBIT:0]  W_7_x251 =  23'd900;
localparam signed [DEBIT:0]  W_7_x252 =  23'd978;
localparam signed [DEBIT:0]  W_7_x253 =  23'd974;
localparam signed [DEBIT:0]  W_7_x254 =  23'd964;
localparam signed [DEBIT:0]  W_7_x255 =  23'd951;
localparam signed [DEBIT:0]  W_7_x256 =  23'd851;
localparam signed [DEBIT:0]  W_7_x257 =  23'd632;
localparam signed [DEBIT:0]  W_7_x258 =  23'd338;
localparam signed [DEBIT:0]  W_7_x259 =  23'd12;
localparam signed [DEBIT:0]  W_7_x260 =  23'd13;
localparam signed [DEBIT:0]  W_7_x261 =  23'd53;
localparam signed [DEBIT:0]  W_7_x262 =  23'd55;
localparam signed [DEBIT:0]  W_7_x263 =  23'd93;
localparam signed [DEBIT:0]  W_7_x264 =  23'd157;
localparam signed [DEBIT:0]  W_7_x265 =  23'd156;
localparam signed [DEBIT:0]  W_7_x266 =  23'd90;
localparam signed [DEBIT:0]  W_7_x267 =  23'd178;
localparam signed [DEBIT:0]  W_7_x268 =  23'd236;
localparam signed [DEBIT:0]  W_7_x269 =  23'd226;
localparam signed [DEBIT:0]  W_7_x270 =  23'd157;
localparam signed [DEBIT:0]  W_7_x271 =  23'd10;
localparam signed [DEBIT:0]  W_7_x272 = - 23'd16;
localparam signed [DEBIT:0]  W_7_x273 = - 23'd44;
localparam signed [DEBIT:0]  W_7_x274 = - 23'd156;
localparam signed [DEBIT:0]  W_7_x275 = - 23'd114;
localparam signed [DEBIT:0]  W_7_x276 =  23'd141;
localparam signed [DEBIT:0]  W_7_x277 =  23'd521;
localparam signed [DEBIT:0]  W_7_x278 =  23'd763;
localparam signed [DEBIT:0]  W_7_x279 =  23'd931;
localparam signed [DEBIT:0]  W_7_x280 =  23'd994;
localparam signed [DEBIT:0]  W_7_x281 =  23'd978;
localparam signed [DEBIT:0]  W_7_x282 =  23'd980;
localparam signed [DEBIT:0]  W_7_x283 =  23'd963;
localparam signed [DEBIT:0]  W_7_x284 =  23'd857;
localparam signed [DEBIT:0]  W_7_x285 =  23'd660;
localparam signed [DEBIT:0]  W_7_x286 =  23'd258;
localparam signed [DEBIT:0]  W_7_x287 = - 23'd72;
localparam signed [DEBIT:0]  W_7_x288 = - 23'd126;
localparam signed [DEBIT:0]  W_7_x289 = - 23'd82;
localparam signed [DEBIT:0]  W_7_x290 = - 23'd59;
localparam signed [DEBIT:0]  W_7_x291 = - 23'd30;
localparam signed [DEBIT:0]  W_7_x292 =  23'd58;
localparam signed [DEBIT:0]  W_7_x293 =  23'd155;
localparam signed [DEBIT:0]  W_7_x294 =  23'd202;
localparam signed [DEBIT:0]  W_7_x295 =  23'd137;
localparam signed [DEBIT:0]  W_7_x296 =  23'd137;
localparam signed [DEBIT:0]  W_7_x297 =  23'd183;
localparam signed [DEBIT:0]  W_7_x298 =  23'd147;
localparam signed [DEBIT:0]  W_7_x299 =  23'd117;
localparam signed [DEBIT:0]  W_7_x300 =  23'd84;
localparam signed [DEBIT:0]  W_7_x301 =  23'd59;
localparam signed [DEBIT:0]  W_7_x302 = - 23'd17;
localparam signed [DEBIT:0]  W_7_x303 =  23'd5;
localparam signed [DEBIT:0]  W_7_x304 =  23'd253;
localparam signed [DEBIT:0]  W_7_x305 =  23'd607;
localparam signed [DEBIT:0]  W_7_x306 =  23'd825;
localparam signed [DEBIT:0]  W_7_x307 =  23'd936;
localparam signed [DEBIT:0]  W_7_x308 =  23'd976;
localparam signed [DEBIT:0]  W_7_x309 =  23'd977;
localparam signed [DEBIT:0]  W_7_x310 =  23'd986;
localparam signed [DEBIT:0]  W_7_x311 =  23'd970;
localparam signed [DEBIT:0]  W_7_x312 =  23'd899;
localparam signed [DEBIT:0]  W_7_x313 =  23'd648;
localparam signed [DEBIT:0]  W_7_x314 =  23'd118;
localparam signed [DEBIT:0]  W_7_x315 = - 23'd190;
localparam signed [DEBIT:0]  W_7_x316 = - 23'd186;
localparam signed [DEBIT:0]  W_7_x317 = - 23'd89;
localparam signed [DEBIT:0]  W_7_x318 = - 23'd2;
localparam signed [DEBIT:0]  W_7_x319 = - 23'd14;
localparam signed [DEBIT:0]  W_7_x320 =  23'd50;
localparam signed [DEBIT:0]  W_7_x321 =  23'd60;
localparam signed [DEBIT:0]  W_7_x322 =  23'd17;
localparam signed [DEBIT:0]  W_7_x323 = - 23'd119;
localparam signed [DEBIT:0]  W_7_x324 =  23'd49;
localparam signed [DEBIT:0]  W_7_x325 =  23'd190;
localparam signed [DEBIT:0]  W_7_x326 =  23'd168;
localparam signed [DEBIT:0]  W_7_x327 =  23'd190;
localparam signed [DEBIT:0]  W_7_x328 =  23'd52;
localparam signed [DEBIT:0]  W_7_x329 = - 23'd22;
localparam signed [DEBIT:0]  W_7_x330 = - 23'd65;
localparam signed [DEBIT:0]  W_7_x331 = - 23'd17;
localparam signed [DEBIT:0]  W_7_x332 =  23'd227;
localparam signed [DEBIT:0]  W_7_x333 =  23'd619;
localparam signed [DEBIT:0]  W_7_x334 =  23'd846;
localparam signed [DEBIT:0]  W_7_x335 =  23'd952;
localparam signed [DEBIT:0]  W_7_x336 =  23'd971;
localparam signed [DEBIT:0]  W_7_x337 =  23'd984;
localparam signed [DEBIT:0]  W_7_x338 =  23'd983;
localparam signed [DEBIT:0]  W_7_x339 =  23'd982;
localparam signed [DEBIT:0]  W_7_x340 =  23'd907;
localparam signed [DEBIT:0]  W_7_x341 =  23'd645;
localparam signed [DEBIT:0]  W_7_x342 =  23'd61;
localparam signed [DEBIT:0]  W_7_x343 = - 23'd235;
localparam signed [DEBIT:0]  W_7_x344 = - 23'd135;
localparam signed [DEBIT:0]  W_7_x345 =  23'd0;
localparam signed [DEBIT:0]  W_7_x346 = - 23'd126;
localparam signed [DEBIT:0]  W_7_x347 = - 23'd266;
localparam signed [DEBIT:0]  W_7_x348 = - 23'd228;
localparam signed [DEBIT:0]  W_7_x349 = - 23'd264;
localparam signed [DEBIT:0]  W_7_x350 = - 23'd410;
localparam signed [DEBIT:0]  W_7_x351 = - 23'd503;
localparam signed [DEBIT:0]  W_7_x352 = - 23'd183;
localparam signed [DEBIT:0]  W_7_x353 =  23'd90;
localparam signed [DEBIT:0]  W_7_x354 =  23'd70;
localparam signed [DEBIT:0]  W_7_x355 =  23'd44;
localparam signed [DEBIT:0]  W_7_x356 = - 23'd10;
localparam signed [DEBIT:0]  W_7_x357 = - 23'd88;
localparam signed [DEBIT:0]  W_7_x358 = - 23'd76;
localparam signed [DEBIT:0]  W_7_x359 =  23'd9;
localparam signed [DEBIT:0]  W_7_x360 =  23'd175;
localparam signed [DEBIT:0]  W_7_x361 =  23'd569;
localparam signed [DEBIT:0]  W_7_x362 =  23'd888;
localparam signed [DEBIT:0]  W_7_x363 =  23'd968;
localparam signed [DEBIT:0]  W_7_x364 =  23'd982;
localparam signed [DEBIT:0]  W_7_x365 =  23'd976;
localparam signed [DEBIT:0]  W_7_x366 =  23'd968;
localparam signed [DEBIT:0]  W_7_x367 =  23'd972;
localparam signed [DEBIT:0]  W_7_x368 =  23'd876;
localparam signed [DEBIT:0]  W_7_x369 =  23'd656;
localparam signed [DEBIT:0]  W_7_x370 =  23'd63;
localparam signed [DEBIT:0]  W_7_x371 = - 23'd266;
localparam signed [DEBIT:0]  W_7_x372 = - 23'd231;
localparam signed [DEBIT:0]  W_7_x373 = - 23'd157;
localparam signed [DEBIT:0]  W_7_x374 = - 23'd302;
localparam signed [DEBIT:0]  W_7_x375 = - 23'd426;
localparam signed [DEBIT:0]  W_7_x376 = - 23'd468;
localparam signed [DEBIT:0]  W_7_x377 = - 23'd525;
localparam signed [DEBIT:0]  W_7_x378 = - 23'd712;
localparam signed [DEBIT:0]  W_7_x379 = - 23'd650;
localparam signed [DEBIT:0]  W_7_x380 = - 23'd255;
localparam signed [DEBIT:0]  W_7_x381 = - 23'd34;
localparam signed [DEBIT:0]  W_7_x382 = - 23'd128;
localparam signed [DEBIT:0]  W_7_x383 = - 23'd166;
localparam signed [DEBIT:0]  W_7_x384 =  23'd6;
localparam signed [DEBIT:0]  W_7_x385 = - 23'd40;
localparam signed [DEBIT:0]  W_7_x386 = - 23'd73;
localparam signed [DEBIT:0]  W_7_x387 =  23'd8;
localparam signed [DEBIT:0]  W_7_x388 =  23'd188;
localparam signed [DEBIT:0]  W_7_x389 =  23'd538;
localparam signed [DEBIT:0]  W_7_x390 =  23'd876;
localparam signed [DEBIT:0]  W_7_x391 =  23'd977;
localparam signed [DEBIT:0]  W_7_x392 =  23'd980;
localparam signed [DEBIT:0]  W_7_x393 =  23'd980;
localparam signed [DEBIT:0]  W_7_x394 =  23'd975;
localparam signed [DEBIT:0]  W_7_x395 =  23'd975;
localparam signed [DEBIT:0]  W_7_x396 =  23'd852;
localparam signed [DEBIT:0]  W_7_x397 =  23'd627;
localparam signed [DEBIT:0]  W_7_x398 =  23'd131;
localparam signed [DEBIT:0]  W_7_x399 = - 23'd293;
localparam signed [DEBIT:0]  W_7_x400 = - 23'd290;
localparam signed [DEBIT:0]  W_7_x401 = - 23'd246;
localparam signed [DEBIT:0]  W_7_x402 = - 23'd360;
localparam signed [DEBIT:0]  W_7_x403 = - 23'd484;
localparam signed [DEBIT:0]  W_7_x404 = - 23'd492;
localparam signed [DEBIT:0]  W_7_x405 = - 23'd543;
localparam signed [DEBIT:0]  W_7_x406 = - 23'd599;
localparam signed [DEBIT:0]  W_7_x407 = - 23'd372;
localparam signed [DEBIT:0]  W_7_x408 = - 23'd112;
localparam signed [DEBIT:0]  W_7_x409 = - 23'd31;
localparam signed [DEBIT:0]  W_7_x410 = - 23'd209;
localparam signed [DEBIT:0]  W_7_x411 =  23'd51;
localparam signed [DEBIT:0]  W_7_x412 =  23'd189;
localparam signed [DEBIT:0]  W_7_x413 =  23'd76;
localparam signed [DEBIT:0]  W_7_x414 =  23'd81;
localparam signed [DEBIT:0]  W_7_x415 =  23'd176;
localparam signed [DEBIT:0]  W_7_x416 =  23'd281;
localparam signed [DEBIT:0]  W_7_x417 =  23'd529;
localparam signed [DEBIT:0]  W_7_x418 =  23'd884;
localparam signed [DEBIT:0]  W_7_x419 =  23'd963;
localparam signed [DEBIT:0]  W_7_x420 =  23'd977;
localparam signed [DEBIT:0]  W_7_x421 =  23'd987;
localparam signed [DEBIT:0]  W_7_x422 =  23'd976;
localparam signed [DEBIT:0]  W_7_x423 =  23'd965;
localparam signed [DEBIT:0]  W_7_x424 =  23'd859;
localparam signed [DEBIT:0]  W_7_x425 =  23'd666;
localparam signed [DEBIT:0]  W_7_x426 =  23'd111;
localparam signed [DEBIT:0]  W_7_x427 = - 23'd225;
localparam signed [DEBIT:0]  W_7_x428 = - 23'd286;
localparam signed [DEBIT:0]  W_7_x429 = - 23'd299;
localparam signed [DEBIT:0]  W_7_x430 = - 23'd294;
localparam signed [DEBIT:0]  W_7_x431 = - 23'd362;
localparam signed [DEBIT:0]  W_7_x432 = - 23'd366;
localparam signed [DEBIT:0]  W_7_x433 = - 23'd330;
localparam signed [DEBIT:0]  W_7_x434 = - 23'd376;
localparam signed [DEBIT:0]  W_7_x435 = - 23'd150;
localparam signed [DEBIT:0]  W_7_x436 = - 23'd13;
localparam signed [DEBIT:0]  W_7_x437 = - 23'd44;
localparam signed [DEBIT:0]  W_7_x438 =  23'd75;
localparam signed [DEBIT:0]  W_7_x439 =  23'd315;
localparam signed [DEBIT:0]  W_7_x440 =  23'd258;
localparam signed [DEBIT:0]  W_7_x441 =  23'd192;
localparam signed [DEBIT:0]  W_7_x442 =  23'd198;
localparam signed [DEBIT:0]  W_7_x443 =  23'd197;
localparam signed [DEBIT:0]  W_7_x444 =  23'd214;
localparam signed [DEBIT:0]  W_7_x445 =  23'd474;
localparam signed [DEBIT:0]  W_7_x446 =  23'd841;
localparam signed [DEBIT:0]  W_7_x447 =  23'd943;
localparam signed [DEBIT:0]  W_7_x448 =  23'd970;
localparam signed [DEBIT:0]  W_7_x449 =  23'd988;
localparam signed [DEBIT:0]  W_7_x450 =  23'd975;
localparam signed [DEBIT:0]  W_7_x451 =  23'd975;
localparam signed [DEBIT:0]  W_7_x452 =  23'd894;
localparam signed [DEBIT:0]  W_7_x453 =  23'd701;
localparam signed [DEBIT:0]  W_7_x454 =  23'd144;
localparam signed [DEBIT:0]  W_7_x455 = - 23'd198;
localparam signed [DEBIT:0]  W_7_x456 = - 23'd229;
localparam signed [DEBIT:0]  W_7_x457 = - 23'd206;
localparam signed [DEBIT:0]  W_7_x458 = - 23'd261;
localparam signed [DEBIT:0]  W_7_x459 = - 23'd271;
localparam signed [DEBIT:0]  W_7_x460 = - 23'd329;
localparam signed [DEBIT:0]  W_7_x461 = - 23'd242;
localparam signed [DEBIT:0]  W_7_x462 = - 23'd248;
localparam signed [DEBIT:0]  W_7_x463 = - 23'd156;
localparam signed [DEBIT:0]  W_7_x464 =  23'd65;
localparam signed [DEBIT:0]  W_7_x465 = - 23'd15;
localparam signed [DEBIT:0]  W_7_x466 =  23'd211;
localparam signed [DEBIT:0]  W_7_x467 =  23'd234;
localparam signed [DEBIT:0]  W_7_x468 =  23'd123;
localparam signed [DEBIT:0]  W_7_x469 =  23'd73;
localparam signed [DEBIT:0]  W_7_x470 =  23'd60;
localparam signed [DEBIT:0]  W_7_x471 =  23'd118;
localparam signed [DEBIT:0]  W_7_x472 =  23'd167;
localparam signed [DEBIT:0]  W_7_x473 =  23'd399;
localparam signed [DEBIT:0]  W_7_x474 =  23'd806;
localparam signed [DEBIT:0]  W_7_x475 =  23'd946;
localparam signed [DEBIT:0]  W_7_x476 =  23'd980;
localparam signed [DEBIT:0]  W_7_x477 =  23'd987;
localparam signed [DEBIT:0]  W_7_x478 =  23'd983;
localparam signed [DEBIT:0]  W_7_x479 =  23'd965;
localparam signed [DEBIT:0]  W_7_x480 =  23'd882;
localparam signed [DEBIT:0]  W_7_x481 =  23'd622;
localparam signed [DEBIT:0]  W_7_x482 =  23'd135;
localparam signed [DEBIT:0]  W_7_x483 = - 23'd167;
localparam signed [DEBIT:0]  W_7_x484 = - 23'd267;
localparam signed [DEBIT:0]  W_7_x485 = - 23'd256;
localparam signed [DEBIT:0]  W_7_x486 = - 23'd203;
localparam signed [DEBIT:0]  W_7_x487 = - 23'd250;
localparam signed [DEBIT:0]  W_7_x488 = - 23'd209;
localparam signed [DEBIT:0]  W_7_x489 = - 23'd142;
localparam signed [DEBIT:0]  W_7_x490 = - 23'd81;
localparam signed [DEBIT:0]  W_7_x491 =  23'd79;
localparam signed [DEBIT:0]  W_7_x492 =  23'd100;
localparam signed [DEBIT:0]  W_7_x493 = - 23'd25;
localparam signed [DEBIT:0]  W_7_x494 =  23'd72;
localparam signed [DEBIT:0]  W_7_x495 =  23'd59;
localparam signed [DEBIT:0]  W_7_x496 = - 23'd121;
localparam signed [DEBIT:0]  W_7_x497 = - 23'd321;
localparam signed [DEBIT:0]  W_7_x498 = - 23'd208;
localparam signed [DEBIT:0]  W_7_x499 = - 23'd53;
localparam signed [DEBIT:0]  W_7_x500 =  23'd144;
localparam signed [DEBIT:0]  W_7_x501 =  23'd451;
localparam signed [DEBIT:0]  W_7_x502 =  23'd832;
localparam signed [DEBIT:0]  W_7_x503 =  23'd961;
localparam signed [DEBIT:0]  W_7_x504 =  23'd975;
localparam signed [DEBIT:0]  W_7_x505 =  23'd982;
localparam signed [DEBIT:0]  W_7_x506 =  23'd986;
localparam signed [DEBIT:0]  W_7_x507 =  23'd963;
localparam signed [DEBIT:0]  W_7_x508 =  23'd845;
localparam signed [DEBIT:0]  W_7_x509 =  23'd545;
localparam signed [DEBIT:0]  W_7_x510 =  23'd69;
localparam signed [DEBIT:0]  W_7_x511 = - 23'd181;
localparam signed [DEBIT:0]  W_7_x512 = - 23'd207;
localparam signed [DEBIT:0]  W_7_x513 = - 23'd197;
localparam signed [DEBIT:0]  W_7_x514 = - 23'd235;
localparam signed [DEBIT:0]  W_7_x515 = - 23'd218;
localparam signed [DEBIT:0]  W_7_x516 =  23'd10;
localparam signed [DEBIT:0]  W_7_x517 =  23'd71;
localparam signed [DEBIT:0]  W_7_x518 =  23'd139;
localparam signed [DEBIT:0]  W_7_x519 =  23'd97;
localparam signed [DEBIT:0]  W_7_x520 = - 23'd125;
localparam signed [DEBIT:0]  W_7_x521 = - 23'd251;
localparam signed [DEBIT:0]  W_7_x522 = - 23'd172;
localparam signed [DEBIT:0]  W_7_x523 = - 23'd127;
localparam signed [DEBIT:0]  W_7_x524 = - 23'd349;
localparam signed [DEBIT:0]  W_7_x525 = - 23'd392;
localparam signed [DEBIT:0]  W_7_x526 = - 23'd388;
localparam signed [DEBIT:0]  W_7_x527 = - 23'd232;
localparam signed [DEBIT:0]  W_7_x528 =  23'd94;
localparam signed [DEBIT:0]  W_7_x529 =  23'd516;
localparam signed [DEBIT:0]  W_7_x530 =  23'd872;
localparam signed [DEBIT:0]  W_7_x531 =  23'd967;
localparam signed [DEBIT:0]  W_7_x532 =  23'd975;
localparam signed [DEBIT:0]  W_7_x533 =  23'd987;
localparam signed [DEBIT:0]  W_7_x534 =  23'd976;
localparam signed [DEBIT:0]  W_7_x535 =  23'd939;
localparam signed [DEBIT:0]  W_7_x536 =  23'd762;
localparam signed [DEBIT:0]  W_7_x537 =  23'd447;
localparam signed [DEBIT:0]  W_7_x538 =  23'd58;
localparam signed [DEBIT:0]  W_7_x539 = - 23'd167;
localparam signed [DEBIT:0]  W_7_x540 = - 23'd212;
localparam signed [DEBIT:0]  W_7_x541 = - 23'd235;
localparam signed [DEBIT:0]  W_7_x542 = - 23'd253;
localparam signed [DEBIT:0]  W_7_x543 = - 23'd152;
localparam signed [DEBIT:0]  W_7_x544 = - 23'd89;
localparam signed [DEBIT:0]  W_7_x545 =  23'd20;
localparam signed [DEBIT:0]  W_7_x546 = - 23'd9;
localparam signed [DEBIT:0]  W_7_x547 = - 23'd60;
localparam signed [DEBIT:0]  W_7_x548 = - 23'd181;
localparam signed [DEBIT:0]  W_7_x549 = - 23'd324;
localparam signed [DEBIT:0]  W_7_x550 = - 23'd265;
localparam signed [DEBIT:0]  W_7_x551 = - 23'd367;
localparam signed [DEBIT:0]  W_7_x552 = - 23'd542;
localparam signed [DEBIT:0]  W_7_x553 = - 23'd558;
localparam signed [DEBIT:0]  W_7_x554 = - 23'd554;
localparam signed [DEBIT:0]  W_7_x555 = - 23'd275;
localparam signed [DEBIT:0]  W_7_x556 =  23'd133;
localparam signed [DEBIT:0]  W_7_x557 =  23'd653;
localparam signed [DEBIT:0]  W_7_x558 =  23'd914;
localparam signed [DEBIT:0]  W_7_x559 =  23'd963;
localparam signed [DEBIT:0]  W_7_x560 =  23'd982;
localparam signed [DEBIT:0]  W_7_x561 =  23'd977;
localparam signed [DEBIT:0]  W_7_x562 =  23'd964;
localparam signed [DEBIT:0]  W_7_x563 =  23'd926;
localparam signed [DEBIT:0]  W_7_x564 =  23'd733;
localparam signed [DEBIT:0]  W_7_x565 =  23'd373;
localparam signed [DEBIT:0]  W_7_x566 =  23'd60;
localparam signed [DEBIT:0]  W_7_x567 = - 23'd201;
localparam signed [DEBIT:0]  W_7_x568 = - 23'd289;
localparam signed [DEBIT:0]  W_7_x569 = - 23'd282;
localparam signed [DEBIT:0]  W_7_x570 = - 23'd254;
localparam signed [DEBIT:0]  W_7_x571 = - 23'd181;
localparam signed [DEBIT:0]  W_7_x572 = - 23'd200;
localparam signed [DEBIT:0]  W_7_x573 = - 23'd101;
localparam signed [DEBIT:0]  W_7_x574 = - 23'd77;
localparam signed [DEBIT:0]  W_7_x575 = - 23'd164;
localparam signed [DEBIT:0]  W_7_x576 = - 23'd256;
localparam signed [DEBIT:0]  W_7_x577 = - 23'd334;
localparam signed [DEBIT:0]  W_7_x578 = - 23'd273;
localparam signed [DEBIT:0]  W_7_x579 = - 23'd404;
localparam signed [DEBIT:0]  W_7_x580 = - 23'd611;
localparam signed [DEBIT:0]  W_7_x581 = - 23'd701;
localparam signed [DEBIT:0]  W_7_x582 = - 23'd497;
localparam signed [DEBIT:0]  W_7_x583 = - 23'd171;
localparam signed [DEBIT:0]  W_7_x584 =  23'd294;
localparam signed [DEBIT:0]  W_7_x585 =  23'd750;
localparam signed [DEBIT:0]  W_7_x586 =  23'd931;
localparam signed [DEBIT:0]  W_7_x587 =  23'd977;
localparam signed [DEBIT:0]  W_7_x588 =  23'd973;
localparam signed [DEBIT:0]  W_7_x589 =  23'd975;
localparam signed [DEBIT:0]  W_7_x590 =  23'd967;
localparam signed [DEBIT:0]  W_7_x591 =  23'd915;
localparam signed [DEBIT:0]  W_7_x592 =  23'd755;
localparam signed [DEBIT:0]  W_7_x593 =  23'd430;
localparam signed [DEBIT:0]  W_7_x594 =  23'd72;
localparam signed [DEBIT:0]  W_7_x595 = - 23'd230;
localparam signed [DEBIT:0]  W_7_x596 = - 23'd444;
localparam signed [DEBIT:0]  W_7_x597 = - 23'd369;
localparam signed [DEBIT:0]  W_7_x598 = - 23'd279;
localparam signed [DEBIT:0]  W_7_x599 = - 23'd235;
localparam signed [DEBIT:0]  W_7_x600 = - 23'd42;
localparam signed [DEBIT:0]  W_7_x601 = - 23'd12;
localparam signed [DEBIT:0]  W_7_x602 = - 23'd26;
localparam signed [DEBIT:0]  W_7_x603 = - 23'd89;
localparam signed [DEBIT:0]  W_7_x604 = - 23'd155;
localparam signed [DEBIT:0]  W_7_x605 = - 23'd216;
localparam signed [DEBIT:0]  W_7_x606 = - 23'd227;
localparam signed [DEBIT:0]  W_7_x607 = - 23'd378;
localparam signed [DEBIT:0]  W_7_x608 = - 23'd577;
localparam signed [DEBIT:0]  W_7_x609 = - 23'd639;
localparam signed [DEBIT:0]  W_7_x610 = - 23'd397;
localparam signed [DEBIT:0]  W_7_x611 = - 23'd46;
localparam signed [DEBIT:0]  W_7_x612 =  23'd475;
localparam signed [DEBIT:0]  W_7_x613 =  23'd762;
localparam signed [DEBIT:0]  W_7_x614 =  23'd941;
localparam signed [DEBIT:0]  W_7_x615 =  23'd979;
localparam signed [DEBIT:0]  W_7_x616 =  23'd977;
localparam signed [DEBIT:0]  W_7_x617 =  23'd974;
localparam signed [DEBIT:0]  W_7_x618 =  23'd975;
localparam signed [DEBIT:0]  W_7_x619 =  23'd932;
localparam signed [DEBIT:0]  W_7_x620 =  23'd829;
localparam signed [DEBIT:0]  W_7_x621 =  23'd580;
localparam signed [DEBIT:0]  W_7_x622 =  23'd299;
localparam signed [DEBIT:0]  W_7_x623 =  23'd3;
localparam signed [DEBIT:0]  W_7_x624 = - 23'd210;
localparam signed [DEBIT:0]  W_7_x625 = - 23'd178;
localparam signed [DEBIT:0]  W_7_x626 = - 23'd99;
localparam signed [DEBIT:0]  W_7_x627 =  23'd7;
localparam signed [DEBIT:0]  W_7_x628 = - 23'd8;
localparam signed [DEBIT:0]  W_7_x629 =  23'd27;
localparam signed [DEBIT:0]  W_7_x630 = - 23'd40;
localparam signed [DEBIT:0]  W_7_x631 = - 23'd6;
localparam signed [DEBIT:0]  W_7_x632 =  23'd43;
localparam signed [DEBIT:0]  W_7_x633 = - 23'd66;
localparam signed [DEBIT:0]  W_7_x634 = - 23'd160;
localparam signed [DEBIT:0]  W_7_x635 = - 23'd347;
localparam signed [DEBIT:0]  W_7_x636 = - 23'd499;
localparam signed [DEBIT:0]  W_7_x637 = - 23'd486;
localparam signed [DEBIT:0]  W_7_x638 = - 23'd207;
localparam signed [DEBIT:0]  W_7_x639 =  23'd212;
localparam signed [DEBIT:0]  W_7_x640 =  23'd611;
localparam signed [DEBIT:0]  W_7_x641 =  23'd835;
localparam signed [DEBIT:0]  W_7_x642 =  23'd947;
localparam signed [DEBIT:0]  W_7_x643 =  23'd972;
localparam signed [DEBIT:0]  W_7_x644 =  23'd988;
localparam signed [DEBIT:0]  W_7_x645 =  23'd982;
localparam signed [DEBIT:0]  W_7_x646 =  23'd977;
localparam signed [DEBIT:0]  W_7_x647 =  23'd958;
localparam signed [DEBIT:0]  W_7_x648 =  23'd894;
localparam signed [DEBIT:0]  W_7_x649 =  23'd786;
localparam signed [DEBIT:0]  W_7_x650 =  23'd594;
localparam signed [DEBIT:0]  W_7_x651 =  23'd393;
localparam signed [DEBIT:0]  W_7_x652 =  23'd251;
localparam signed [DEBIT:0]  W_7_x653 =  23'd116;
localparam signed [DEBIT:0]  W_7_x654 =  23'd28;
localparam signed [DEBIT:0]  W_7_x655 =  23'd52;
localparam signed [DEBIT:0]  W_7_x656 =  23'd11;
localparam signed [DEBIT:0]  W_7_x657 =  23'd73;
localparam signed [DEBIT:0]  W_7_x658 =  23'd20;
localparam signed [DEBIT:0]  W_7_x659 =  23'd62;
localparam signed [DEBIT:0]  W_7_x660 =  23'd97;
localparam signed [DEBIT:0]  W_7_x661 =  23'd57;
localparam signed [DEBIT:0]  W_7_x662 = - 23'd21;
localparam signed [DEBIT:0]  W_7_x663 = - 23'd162;
localparam signed [DEBIT:0]  W_7_x664 = - 23'd173;
localparam signed [DEBIT:0]  W_7_x665 = - 23'd99;
localparam signed [DEBIT:0]  W_7_x666 =  23'd146;
localparam signed [DEBIT:0]  W_7_x667 =  23'd459;
localparam signed [DEBIT:0]  W_7_x668 =  23'd737;
localparam signed [DEBIT:0]  W_7_x669 =  23'd905;
localparam signed [DEBIT:0]  W_7_x670 =  23'd961;
localparam signed [DEBIT:0]  W_7_x671 =  23'd969;
localparam signed [DEBIT:0]  W_7_x672 =  23'd978;
localparam signed [DEBIT:0]  W_7_x673 =  23'd979;
localparam signed [DEBIT:0]  W_7_x674 =  23'd976;
localparam signed [DEBIT:0]  W_7_x675 =  23'd967;
localparam signed [DEBIT:0]  W_7_x676 =  23'd946;
localparam signed [DEBIT:0]  W_7_x677 =  23'd907;
localparam signed [DEBIT:0]  W_7_x678 =  23'd857;
localparam signed [DEBIT:0]  W_7_x679 =  23'd784;
localparam signed [DEBIT:0]  W_7_x680 =  23'd680;
localparam signed [DEBIT:0]  W_7_x681 =  23'd541;
localparam signed [DEBIT:0]  W_7_x682 =  23'd372;
localparam signed [DEBIT:0]  W_7_x683 =  23'd326;
localparam signed [DEBIT:0]  W_7_x684 =  23'd307;
localparam signed [DEBIT:0]  W_7_x685 =  23'd326;
localparam signed [DEBIT:0]  W_7_x686 =  23'd335;
localparam signed [DEBIT:0]  W_7_x687 =  23'd438;
localparam signed [DEBIT:0]  W_7_x688 =  23'd348;
localparam signed [DEBIT:0]  W_7_x689 =  23'd282;
localparam signed [DEBIT:0]  W_7_x690 =  23'd349;
localparam signed [DEBIT:0]  W_7_x691 =  23'd283;
localparam signed [DEBIT:0]  W_7_x692 =  23'd356;
localparam signed [DEBIT:0]  W_7_x693 =  23'd387;
localparam signed [DEBIT:0]  W_7_x694 =  23'd471;
localparam signed [DEBIT:0]  W_7_x695 =  23'd652;
localparam signed [DEBIT:0]  W_7_x696 =  23'd825;
localparam signed [DEBIT:0]  W_7_x697 =  23'd939;
localparam signed [DEBIT:0]  W_7_x698 =  23'd961;
localparam signed [DEBIT:0]  W_7_x699 =  23'd983;
localparam signed [DEBIT:0]  W_7_x700 =  23'd976;
localparam signed [DEBIT:0]  W_7_x701 =  23'd975;
localparam signed [DEBIT:0]  W_7_x702 =  23'd974;
localparam signed [DEBIT:0]  W_7_x703 =  23'd978;
localparam signed [DEBIT:0]  W_7_x704 =  23'd981;
localparam signed [DEBIT:0]  W_7_x705 =  23'd977;
localparam signed [DEBIT:0]  W_7_x706 =  23'd961;
localparam signed [DEBIT:0]  W_7_x707 =  23'd929;
localparam signed [DEBIT:0]  W_7_x708 =  23'd940;
localparam signed [DEBIT:0]  W_7_x709 =  23'd865;
localparam signed [DEBIT:0]  W_7_x710 =  23'd762;
localparam signed [DEBIT:0]  W_7_x711 =  23'd698;
localparam signed [DEBIT:0]  W_7_x712 =  23'd643;
localparam signed [DEBIT:0]  W_7_x713 =  23'd618;
localparam signed [DEBIT:0]  W_7_x714 =  23'd637;
localparam signed [DEBIT:0]  W_7_x715 =  23'd760;
localparam signed [DEBIT:0]  W_7_x716 =  23'd769;
localparam signed [DEBIT:0]  W_7_x717 =  23'd759;
localparam signed [DEBIT:0]  W_7_x718 =  23'd807;
localparam signed [DEBIT:0]  W_7_x719 =  23'd770;
localparam signed [DEBIT:0]  W_7_x720 =  23'd746;
localparam signed [DEBIT:0]  W_7_x721 =  23'd685;
localparam signed [DEBIT:0]  W_7_x722 =  23'd740;
localparam signed [DEBIT:0]  W_7_x723 =  23'd835;
localparam signed [DEBIT:0]  W_7_x724 =  23'd923;
localparam signed [DEBIT:0]  W_7_x725 =  23'd975;
localparam signed [DEBIT:0]  W_7_x726 =  23'd968;
localparam signed [DEBIT:0]  W_7_x727 =  23'd970;
localparam signed [DEBIT:0]  W_7_x728 =  23'd979;
localparam signed [DEBIT:0]  W_7_x729 =  23'd970;
localparam signed [DEBIT:0]  W_7_x730 =  23'd976;
localparam signed [DEBIT:0]  W_7_x731 =  23'd977;
localparam signed [DEBIT:0]  W_7_x732 =  23'd984;
localparam signed [DEBIT:0]  W_7_x733 =  23'd978;
localparam signed [DEBIT:0]  W_7_x734 =  23'd972;
localparam signed [DEBIT:0]  W_7_x735 =  23'd964;
localparam signed [DEBIT:0]  W_7_x736 =  23'd973;
localparam signed [DEBIT:0]  W_7_x737 =  23'd962;
localparam signed [DEBIT:0]  W_7_x738 =  23'd914;
localparam signed [DEBIT:0]  W_7_x739 =  23'd853;
localparam signed [DEBIT:0]  W_7_x740 =  23'd794;
localparam signed [DEBIT:0]  W_7_x741 =  23'd756;
localparam signed [DEBIT:0]  W_7_x742 =  23'd782;
localparam signed [DEBIT:0]  W_7_x743 =  23'd815;
localparam signed [DEBIT:0]  W_7_x744 =  23'd887;
localparam signed [DEBIT:0]  W_7_x745 =  23'd889;
localparam signed [DEBIT:0]  W_7_x746 =  23'd901;
localparam signed [DEBIT:0]  W_7_x747 =  23'd898;
localparam signed [DEBIT:0]  W_7_x748 =  23'd896;
localparam signed [DEBIT:0]  W_7_x749 =  23'd851;
localparam signed [DEBIT:0]  W_7_x750 =  23'd893;
localparam signed [DEBIT:0]  W_7_x751 =  23'd934;
localparam signed [DEBIT:0]  W_7_x752 =  23'd970;
localparam signed [DEBIT:0]  W_7_x753 =  23'd985;
localparam signed [DEBIT:0]  W_7_x754 =  23'd979;
localparam signed [DEBIT:0]  W_7_x755 =  23'd987;
localparam signed [DEBIT:0]  W_7_x756 =  23'd969;
localparam signed [DEBIT:0]  W_7_x757 =  23'd987;
localparam signed [DEBIT:0]  W_7_x758 =  23'd974;
localparam signed [DEBIT:0]  W_7_x759 =  23'd981;
localparam signed [DEBIT:0]  W_7_x760 =  23'd973;
localparam signed [DEBIT:0]  W_7_x761 =  23'd973;
localparam signed [DEBIT:0]  W_7_x762 =  23'd974;
localparam signed [DEBIT:0]  W_7_x763 =  23'd976;
localparam signed [DEBIT:0]  W_7_x764 =  23'd982;
localparam signed [DEBIT:0]  W_7_x765 =  23'd974;
localparam signed [DEBIT:0]  W_7_x766 =  23'd979;
localparam signed [DEBIT:0]  W_7_x767 =  23'd973;
localparam signed [DEBIT:0]  W_7_x768 =  23'd970;
localparam signed [DEBIT:0]  W_7_x769 =  23'd969;
localparam signed [DEBIT:0]  W_7_x770 =  23'd985;
localparam signed [DEBIT:0]  W_7_x771 =  23'd983;
localparam signed [DEBIT:0]  W_7_x772 =  23'd971;
localparam signed [DEBIT:0]  W_7_x773 =  23'd987;
localparam signed [DEBIT:0]  W_7_x774 =  23'd990;
localparam signed [DEBIT:0]  W_7_x775 =  23'd974;
localparam signed [DEBIT:0]  W_7_x776 =  23'd969;
localparam signed [DEBIT:0]  W_7_x777 =  23'd970;
localparam signed [DEBIT:0]  W_7_x778 =  23'd969;
localparam signed [DEBIT:0]  W_7_x779 =  23'd973;
localparam signed [DEBIT:0]  W_7_x780 =  23'd977;
localparam signed [DEBIT:0]  W_7_x781 =  23'd984;
localparam signed [DEBIT:0]  W_7_x782 =  23'd984;
localparam signed [DEBIT:0]  W_7_x783 =  23'd990;
localparam signed [DEBIT:0]  W_7_x784 =  23'd975;
localparam signed [DEBIT:0]  W_8_x1 =  23'd941;
localparam signed [DEBIT:0]  W_8_x2 =  23'd943;
localparam signed [DEBIT:0]  W_8_x3 =  23'd944;
localparam signed [DEBIT:0]  W_8_x4 =  23'd939;
localparam signed [DEBIT:0]  W_8_x5 =  23'd940;
localparam signed [DEBIT:0]  W_8_x6 =  23'd952;
localparam signed [DEBIT:0]  W_8_x7 =  23'd942;
localparam signed [DEBIT:0]  W_8_x8 =  23'd943;
localparam signed [DEBIT:0]  W_8_x9 =  23'd942;
localparam signed [DEBIT:0]  W_8_x10 =  23'd939;
localparam signed [DEBIT:0]  W_8_x11 =  23'd944;
localparam signed [DEBIT:0]  W_8_x12 =  23'd940;
localparam signed [DEBIT:0]  W_8_x13 =  23'd941;
localparam signed [DEBIT:0]  W_8_x14 =  23'd936;
localparam signed [DEBIT:0]  W_8_x15 =  23'd934;
localparam signed [DEBIT:0]  W_8_x16 =  23'd941;
localparam signed [DEBIT:0]  W_8_x17 =  23'd940;
localparam signed [DEBIT:0]  W_8_x18 =  23'd946;
localparam signed [DEBIT:0]  W_8_x19 =  23'd927;
localparam signed [DEBIT:0]  W_8_x20 =  23'd946;
localparam signed [DEBIT:0]  W_8_x21 =  23'd930;
localparam signed [DEBIT:0]  W_8_x22 =  23'd942;
localparam signed [DEBIT:0]  W_8_x23 =  23'd944;
localparam signed [DEBIT:0]  W_8_x24 =  23'd939;
localparam signed [DEBIT:0]  W_8_x25 =  23'd947;
localparam signed [DEBIT:0]  W_8_x26 =  23'd936;
localparam signed [DEBIT:0]  W_8_x27 =  23'd941;
localparam signed [DEBIT:0]  W_8_x28 =  23'd933;
localparam signed [DEBIT:0]  W_8_x29 =  23'd946;
localparam signed [DEBIT:0]  W_8_x30 =  23'd939;
localparam signed [DEBIT:0]  W_8_x31 =  23'd943;
localparam signed [DEBIT:0]  W_8_x32 =  23'd931;
localparam signed [DEBIT:0]  W_8_x33 =  23'd948;
localparam signed [DEBIT:0]  W_8_x34 =  23'd938;
localparam signed [DEBIT:0]  W_8_x35 =  23'd941;
localparam signed [DEBIT:0]  W_8_x36 =  23'd930;
localparam signed [DEBIT:0]  W_8_x37 =  23'd943;
localparam signed [DEBIT:0]  W_8_x38 =  23'd921;
localparam signed [DEBIT:0]  W_8_x39 =  23'd913;
localparam signed [DEBIT:0]  W_8_x40 =  23'd914;
localparam signed [DEBIT:0]  W_8_x41 =  23'd916;
localparam signed [DEBIT:0]  W_8_x42 =  23'd920;
localparam signed [DEBIT:0]  W_8_x43 =  23'd904;
localparam signed [DEBIT:0]  W_8_x44 =  23'd915;
localparam signed [DEBIT:0]  W_8_x45 =  23'd902;
localparam signed [DEBIT:0]  W_8_x46 =  23'd921;
localparam signed [DEBIT:0]  W_8_x47 =  23'd931;
localparam signed [DEBIT:0]  W_8_x48 =  23'd923;
localparam signed [DEBIT:0]  W_8_x49 =  23'd937;
localparam signed [DEBIT:0]  W_8_x50 =  23'd942;
localparam signed [DEBIT:0]  W_8_x51 =  23'd953;
localparam signed [DEBIT:0]  W_8_x52 =  23'd933;
localparam signed [DEBIT:0]  W_8_x53 =  23'd942;
localparam signed [DEBIT:0]  W_8_x54 =  23'd938;
localparam signed [DEBIT:0]  W_8_x55 =  23'd937;
localparam signed [DEBIT:0]  W_8_x56 =  23'd946;
localparam signed [DEBIT:0]  W_8_x57 =  23'd946;
localparam signed [DEBIT:0]  W_8_x58 =  23'd945;
localparam signed [DEBIT:0]  W_8_x59 =  23'd942;
localparam signed [DEBIT:0]  W_8_x60 =  23'd938;
localparam signed [DEBIT:0]  W_8_x61 =  23'd932;
localparam signed [DEBIT:0]  W_8_x62 =  23'd943;
localparam signed [DEBIT:0]  W_8_x63 =  23'd934;
localparam signed [DEBIT:0]  W_8_x64 =  23'd920;
localparam signed [DEBIT:0]  W_8_x65 =  23'd880;
localparam signed [DEBIT:0]  W_8_x66 =  23'd841;
localparam signed [DEBIT:0]  W_8_x67 =  23'd823;
localparam signed [DEBIT:0]  W_8_x68 =  23'd812;
localparam signed [DEBIT:0]  W_8_x69 =  23'd774;
localparam signed [DEBIT:0]  W_8_x70 =  23'd746;
localparam signed [DEBIT:0]  W_8_x71 =  23'd697;
localparam signed [DEBIT:0]  W_8_x72 =  23'd687;
localparam signed [DEBIT:0]  W_8_x73 =  23'd684;
localparam signed [DEBIT:0]  W_8_x74 =  23'd733;
localparam signed [DEBIT:0]  W_8_x75 =  23'd768;
localparam signed [DEBIT:0]  W_8_x76 =  23'd781;
localparam signed [DEBIT:0]  W_8_x77 =  23'd881;
localparam signed [DEBIT:0]  W_8_x78 =  23'd919;
localparam signed [DEBIT:0]  W_8_x79 =  23'd936;
localparam signed [DEBIT:0]  W_8_x80 =  23'd931;
localparam signed [DEBIT:0]  W_8_x81 =  23'd945;
localparam signed [DEBIT:0]  W_8_x82 =  23'd933;
localparam signed [DEBIT:0]  W_8_x83 =  23'd937;
localparam signed [DEBIT:0]  W_8_x84 =  23'd938;
localparam signed [DEBIT:0]  W_8_x85 =  23'd944;
localparam signed [DEBIT:0]  W_8_x86 =  23'd936;
localparam signed [DEBIT:0]  W_8_x87 =  23'd938;
localparam signed [DEBIT:0]  W_8_x88 =  23'd945;
localparam signed [DEBIT:0]  W_8_x89 =  23'd937;
localparam signed [DEBIT:0]  W_8_x90 =  23'd911;
localparam signed [DEBIT:0]  W_8_x91 =  23'd862;
localparam signed [DEBIT:0]  W_8_x92 =  23'd768;
localparam signed [DEBIT:0]  W_8_x93 =  23'd674;
localparam signed [DEBIT:0]  W_8_x94 =  23'd597;
localparam signed [DEBIT:0]  W_8_x95 =  23'd506;
localparam signed [DEBIT:0]  W_8_x96 =  23'd378;
localparam signed [DEBIT:0]  W_8_x97 =  23'd293;
localparam signed [DEBIT:0]  W_8_x98 =  23'd244;
localparam signed [DEBIT:0]  W_8_x99 =  23'd150;
localparam signed [DEBIT:0]  W_8_x100 =  23'd99;
localparam signed [DEBIT:0]  W_8_x101 =  23'd80;
localparam signed [DEBIT:0]  W_8_x102 =  23'd119;
localparam signed [DEBIT:0]  W_8_x103 =  23'd210;
localparam signed [DEBIT:0]  W_8_x104 =  23'd338;
localparam signed [DEBIT:0]  W_8_x105 =  23'd548;
localparam signed [DEBIT:0]  W_8_x106 =  23'd705;
localparam signed [DEBIT:0]  W_8_x107 =  23'd825;
localparam signed [DEBIT:0]  W_8_x108 =  23'd892;
localparam signed [DEBIT:0]  W_8_x109 =  23'd921;
localparam signed [DEBIT:0]  W_8_x110 =  23'd927;
localparam signed [DEBIT:0]  W_8_x111 =  23'd944;
localparam signed [DEBIT:0]  W_8_x112 =  23'd933;
localparam signed [DEBIT:0]  W_8_x113 =  23'd931;
localparam signed [DEBIT:0]  W_8_x114 =  23'd942;
localparam signed [DEBIT:0]  W_8_x115 =  23'd945;
localparam signed [DEBIT:0]  W_8_x116 =  23'd933;
localparam signed [DEBIT:0]  W_8_x117 =  23'd916;
localparam signed [DEBIT:0]  W_8_x118 =  23'd825;
localparam signed [DEBIT:0]  W_8_x119 =  23'd698;
localparam signed [DEBIT:0]  W_8_x120 =  23'd525;
localparam signed [DEBIT:0]  W_8_x121 =  23'd309;
localparam signed [DEBIT:0]  W_8_x122 =  23'd103;
localparam signed [DEBIT:0]  W_8_x123 =  23'd28;
localparam signed [DEBIT:0]  W_8_x124 = - 23'd40;
localparam signed [DEBIT:0]  W_8_x125 = - 23'd93;
localparam signed [DEBIT:0]  W_8_x126 = - 23'd25;
localparam signed [DEBIT:0]  W_8_x127 =  23'd1;
localparam signed [DEBIT:0]  W_8_x128 = - 23'd41;
localparam signed [DEBIT:0]  W_8_x129 = - 23'd178;
localparam signed [DEBIT:0]  W_8_x130 = - 23'd324;
localparam signed [DEBIT:0]  W_8_x131 = - 23'd278;
localparam signed [DEBIT:0]  W_8_x132 = - 23'd159;
localparam signed [DEBIT:0]  W_8_x133 = - 23'd25;
localparam signed [DEBIT:0]  W_8_x134 =  23'd168;
localparam signed [DEBIT:0]  W_8_x135 =  23'd369;
localparam signed [DEBIT:0]  W_8_x136 =  23'd634;
localparam signed [DEBIT:0]  W_8_x137 =  23'd833;
localparam signed [DEBIT:0]  W_8_x138 =  23'd901;
localparam signed [DEBIT:0]  W_8_x139 =  23'd933;
localparam signed [DEBIT:0]  W_8_x140 =  23'd942;
localparam signed [DEBIT:0]  W_8_x141 =  23'd941;
localparam signed [DEBIT:0]  W_8_x142 =  23'd936;
localparam signed [DEBIT:0]  W_8_x143 =  23'd942;
localparam signed [DEBIT:0]  W_8_x144 =  23'd929;
localparam signed [DEBIT:0]  W_8_x145 =  23'd844;
localparam signed [DEBIT:0]  W_8_x146 =  23'd594;
localparam signed [DEBIT:0]  W_8_x147 =  23'd277;
localparam signed [DEBIT:0]  W_8_x148 = - 23'd41;
localparam signed [DEBIT:0]  W_8_x149 = - 23'd248;
localparam signed [DEBIT:0]  W_8_x150 = - 23'd287;
localparam signed [DEBIT:0]  W_8_x151 = - 23'd310;
localparam signed [DEBIT:0]  W_8_x152 = - 23'd109;
localparam signed [DEBIT:0]  W_8_x153 =  23'd73;
localparam signed [DEBIT:0]  W_8_x154 =  23'd101;
localparam signed [DEBIT:0]  W_8_x155 =  23'd226;
localparam signed [DEBIT:0]  W_8_x156 =  23'd163;
localparam signed [DEBIT:0]  W_8_x157 =  23'd129;
localparam signed [DEBIT:0]  W_8_x158 =  23'd214;
localparam signed [DEBIT:0]  W_8_x159 =  23'd177;
localparam signed [DEBIT:0]  W_8_x160 =  23'd113;
localparam signed [DEBIT:0]  W_8_x161 = - 23'd149;
localparam signed [DEBIT:0]  W_8_x162 = - 23'd249;
localparam signed [DEBIT:0]  W_8_x163 = - 23'd68;
localparam signed [DEBIT:0]  W_8_x164 =  23'd147;
localparam signed [DEBIT:0]  W_8_x165 =  23'd442;
localparam signed [DEBIT:0]  W_8_x166 =  23'd772;
localparam signed [DEBIT:0]  W_8_x167 =  23'd916;
localparam signed [DEBIT:0]  W_8_x168 =  23'd942;
localparam signed [DEBIT:0]  W_8_x169 =  23'd936;
localparam signed [DEBIT:0]  W_8_x170 =  23'd941;
localparam signed [DEBIT:0]  W_8_x171 =  23'd929;
localparam signed [DEBIT:0]  W_8_x172 =  23'd820;
localparam signed [DEBIT:0]  W_8_x173 =  23'd654;
localparam signed [DEBIT:0]  W_8_x174 =  23'd342;
localparam signed [DEBIT:0]  W_8_x175 = - 23'd23;
localparam signed [DEBIT:0]  W_8_x176 = - 23'd275;
localparam signed [DEBIT:0]  W_8_x177 = - 23'd270;
localparam signed [DEBIT:0]  W_8_x178 = - 23'd267;
localparam signed [DEBIT:0]  W_8_x179 = - 23'd199;
localparam signed [DEBIT:0]  W_8_x180 = - 23'd5;
localparam signed [DEBIT:0]  W_8_x181 =  23'd70;
localparam signed [DEBIT:0]  W_8_x182 =  23'd38;
localparam signed [DEBIT:0]  W_8_x183 =  23'd149;
localparam signed [DEBIT:0]  W_8_x184 =  23'd183;
localparam signed [DEBIT:0]  W_8_x185 =  23'd133;
localparam signed [DEBIT:0]  W_8_x186 =  23'd164;
localparam signed [DEBIT:0]  W_8_x187 =  23'd52;
localparam signed [DEBIT:0]  W_8_x188 =  23'd72;
localparam signed [DEBIT:0]  W_8_x189 = - 23'd132;
localparam signed [DEBIT:0]  W_8_x190 = - 23'd189;
localparam signed [DEBIT:0]  W_8_x191 = - 23'd169;
localparam signed [DEBIT:0]  W_8_x192 = - 23'd18;
localparam signed [DEBIT:0]  W_8_x193 =  23'd180;
localparam signed [DEBIT:0]  W_8_x194 =  23'd546;
localparam signed [DEBIT:0]  W_8_x195 =  23'd834;
localparam signed [DEBIT:0]  W_8_x196 =  23'd937;
localparam signed [DEBIT:0]  W_8_x197 =  23'd943;
localparam signed [DEBIT:0]  W_8_x198 =  23'd930;
localparam signed [DEBIT:0]  W_8_x199 =  23'd900;
localparam signed [DEBIT:0]  W_8_x200 =  23'd703;
localparam signed [DEBIT:0]  W_8_x201 =  23'd456;
localparam signed [DEBIT:0]  W_8_x202 =  23'd147;
localparam signed [DEBIT:0]  W_8_x203 = - 23'd121;
localparam signed [DEBIT:0]  W_8_x204 = - 23'd95;
localparam signed [DEBIT:0]  W_8_x205 =  23'd51;
localparam signed [DEBIT:0]  W_8_x206 =  23'd19;
localparam signed [DEBIT:0]  W_8_x207 =  23'd50;
localparam signed [DEBIT:0]  W_8_x208 =  23'd11;
localparam signed [DEBIT:0]  W_8_x209 = - 23'd12;
localparam signed [DEBIT:0]  W_8_x210 = - 23'd91;
localparam signed [DEBIT:0]  W_8_x211 = - 23'd128;
localparam signed [DEBIT:0]  W_8_x212 = - 23'd34;
localparam signed [DEBIT:0]  W_8_x213 = - 23'd14;
localparam signed [DEBIT:0]  W_8_x214 = - 23'd164;
localparam signed [DEBIT:0]  W_8_x215 = - 23'd34;
localparam signed [DEBIT:0]  W_8_x216 = - 23'd8;
localparam signed [DEBIT:0]  W_8_x217 =  23'd45;
localparam signed [DEBIT:0]  W_8_x218 =  23'd22;
localparam signed [DEBIT:0]  W_8_x219 = - 23'd113;
localparam signed [DEBIT:0]  W_8_x220 =  23'd48;
localparam signed [DEBIT:0]  W_8_x221 =  23'd217;
localparam signed [DEBIT:0]  W_8_x222 =  23'd443;
localparam signed [DEBIT:0]  W_8_x223 =  23'd790;
localparam signed [DEBIT:0]  W_8_x224 =  23'd941;
localparam signed [DEBIT:0]  W_8_x225 =  23'd929;
localparam signed [DEBIT:0]  W_8_x226 =  23'd869;
localparam signed [DEBIT:0]  W_8_x227 =  23'd780;
localparam signed [DEBIT:0]  W_8_x228 =  23'd508;
localparam signed [DEBIT:0]  W_8_x229 =  23'd185;
localparam signed [DEBIT:0]  W_8_x230 = - 23'd69;
localparam signed [DEBIT:0]  W_8_x231 = - 23'd160;
localparam signed [DEBIT:0]  W_8_x232 =  23'd62;
localparam signed [DEBIT:0]  W_8_x233 =  23'd82;
localparam signed [DEBIT:0]  W_8_x234 =  23'd149;
localparam signed [DEBIT:0]  W_8_x235 =  23'd54;
localparam signed [DEBIT:0]  W_8_x236 = - 23'd59;
localparam signed [DEBIT:0]  W_8_x237 =  23'd7;
localparam signed [DEBIT:0]  W_8_x238 = - 23'd65;
localparam signed [DEBIT:0]  W_8_x239 = - 23'd234;
localparam signed [DEBIT:0]  W_8_x240 = - 23'd139;
localparam signed [DEBIT:0]  W_8_x241 =  23'd4;
localparam signed [DEBIT:0]  W_8_x242 = - 23'd154;
localparam signed [DEBIT:0]  W_8_x243 = - 23'd83;
localparam signed [DEBIT:0]  W_8_x244 =  23'd20;
localparam signed [DEBIT:0]  W_8_x245 =  23'd24;
localparam signed [DEBIT:0]  W_8_x246 = - 23'd31;
localparam signed [DEBIT:0]  W_8_x247 =  23'd0;
localparam signed [DEBIT:0]  W_8_x248 =  23'd190;
localparam signed [DEBIT:0]  W_8_x249 =  23'd395;
localparam signed [DEBIT:0]  W_8_x250 =  23'd481;
localparam signed [DEBIT:0]  W_8_x251 =  23'd798;
localparam signed [DEBIT:0]  W_8_x252 =  23'd939;
localparam signed [DEBIT:0]  W_8_x253 =  23'd939;
localparam signed [DEBIT:0]  W_8_x254 =  23'd863;
localparam signed [DEBIT:0]  W_8_x255 =  23'd709;
localparam signed [DEBIT:0]  W_8_x256 =  23'd407;
localparam signed [DEBIT:0]  W_8_x257 =  23'd75;
localparam signed [DEBIT:0]  W_8_x258 = - 23'd135;
localparam signed [DEBIT:0]  W_8_x259 = - 23'd147;
localparam signed [DEBIT:0]  W_8_x260 =  23'd59;
localparam signed [DEBIT:0]  W_8_x261 =  23'd90;
localparam signed [DEBIT:0]  W_8_x262 =  23'd114;
localparam signed [DEBIT:0]  W_8_x263 =  23'd66;
localparam signed [DEBIT:0]  W_8_x264 =  23'd27;
localparam signed [DEBIT:0]  W_8_x265 =  23'd33;
localparam signed [DEBIT:0]  W_8_x266 = - 23'd137;
localparam signed [DEBIT:0]  W_8_x267 = - 23'd384;
localparam signed [DEBIT:0]  W_8_x268 = - 23'd458;
localparam signed [DEBIT:0]  W_8_x269 = - 23'd271;
localparam signed [DEBIT:0]  W_8_x270 = - 23'd99;
localparam signed [DEBIT:0]  W_8_x271 = - 23'd74;
localparam signed [DEBIT:0]  W_8_x272 = - 23'd54;
localparam signed [DEBIT:0]  W_8_x273 =  23'd53;
localparam signed [DEBIT:0]  W_8_x274 =  23'd50;
localparam signed [DEBIT:0]  W_8_x275 =  23'd99;
localparam signed [DEBIT:0]  W_8_x276 =  23'd274;
localparam signed [DEBIT:0]  W_8_x277 =  23'd446;
localparam signed [DEBIT:0]  W_8_x278 =  23'd512;
localparam signed [DEBIT:0]  W_8_x279 =  23'd790;
localparam signed [DEBIT:0]  W_8_x280 =  23'd938;
localparam signed [DEBIT:0]  W_8_x281 =  23'd948;
localparam signed [DEBIT:0]  W_8_x282 =  23'd878;
localparam signed [DEBIT:0]  W_8_x283 =  23'd707;
localparam signed [DEBIT:0]  W_8_x284 =  23'd428;
localparam signed [DEBIT:0]  W_8_x285 =  23'd145;
localparam signed [DEBIT:0]  W_8_x286 = - 23'd60;
localparam signed [DEBIT:0]  W_8_x287 = - 23'd14;
localparam signed [DEBIT:0]  W_8_x288 =  23'd141;
localparam signed [DEBIT:0]  W_8_x289 =  23'd170;
localparam signed [DEBIT:0]  W_8_x290 =  23'd134;
localparam signed [DEBIT:0]  W_8_x291 =  23'd158;
localparam signed [DEBIT:0]  W_8_x292 =  23'd71;
localparam signed [DEBIT:0]  W_8_x293 =  23'd208;
localparam signed [DEBIT:0]  W_8_x294 = - 23'd59;
localparam signed [DEBIT:0]  W_8_x295 = - 23'd441;
localparam signed [DEBIT:0]  W_8_x296 = - 23'd534;
localparam signed [DEBIT:0]  W_8_x297 = - 23'd432;
localparam signed [DEBIT:0]  W_8_x298 = - 23'd196;
localparam signed [DEBIT:0]  W_8_x299 = - 23'd110;
localparam signed [DEBIT:0]  W_8_x300 =  23'd51;
localparam signed [DEBIT:0]  W_8_x301 =  23'd40;
localparam signed [DEBIT:0]  W_8_x302 =  23'd182;
localparam signed [DEBIT:0]  W_8_x303 =  23'd223;
localparam signed [DEBIT:0]  W_8_x304 =  23'd399;
localparam signed [DEBIT:0]  W_8_x305 =  23'd583;
localparam signed [DEBIT:0]  W_8_x306 =  23'd671;
localparam signed [DEBIT:0]  W_8_x307 =  23'd853;
localparam signed [DEBIT:0]  W_8_x308 =  23'd937;
localparam signed [DEBIT:0]  W_8_x309 =  23'd935;
localparam signed [DEBIT:0]  W_8_x310 =  23'd896;
localparam signed [DEBIT:0]  W_8_x311 =  23'd752;
localparam signed [DEBIT:0]  W_8_x312 =  23'd497;
localparam signed [DEBIT:0]  W_8_x313 =  23'd258;
localparam signed [DEBIT:0]  W_8_x314 =  23'd45;
localparam signed [DEBIT:0]  W_8_x315 = - 23'd29;
localparam signed [DEBIT:0]  W_8_x316 =  23'd165;
localparam signed [DEBIT:0]  W_8_x317 =  23'd281;
localparam signed [DEBIT:0]  W_8_x318 =  23'd223;
localparam signed [DEBIT:0]  W_8_x319 =  23'd200;
localparam signed [DEBIT:0]  W_8_x320 =  23'd178;
localparam signed [DEBIT:0]  W_8_x321 =  23'd372;
localparam signed [DEBIT:0]  W_8_x322 =  23'd295;
localparam signed [DEBIT:0]  W_8_x323 = - 23'd60;
localparam signed [DEBIT:0]  W_8_x324 = - 23'd95;
localparam signed [DEBIT:0]  W_8_x325 = - 23'd226;
localparam signed [DEBIT:0]  W_8_x326 = - 23'd61;
localparam signed [DEBIT:0]  W_8_x327 =  23'd45;
localparam signed [DEBIT:0]  W_8_x328 =  23'd75;
localparam signed [DEBIT:0]  W_8_x329 =  23'd67;
localparam signed [DEBIT:0]  W_8_x330 =  23'd88;
localparam signed [DEBIT:0]  W_8_x331 =  23'd179;
localparam signed [DEBIT:0]  W_8_x332 =  23'd325;
localparam signed [DEBIT:0]  W_8_x333 =  23'd719;
localparam signed [DEBIT:0]  W_8_x334 =  23'd849;
localparam signed [DEBIT:0]  W_8_x335 =  23'd881;
localparam signed [DEBIT:0]  W_8_x336 =  23'd941;
localparam signed [DEBIT:0]  W_8_x337 =  23'd936;
localparam signed [DEBIT:0]  W_8_x338 =  23'd921;
localparam signed [DEBIT:0]  W_8_x339 =  23'd818;
localparam signed [DEBIT:0]  W_8_x340 =  23'd623;
localparam signed [DEBIT:0]  W_8_x341 =  23'd356;
localparam signed [DEBIT:0]  W_8_x342 =  23'd87;
localparam signed [DEBIT:0]  W_8_x343 = - 23'd30;
localparam signed [DEBIT:0]  W_8_x344 =  23'd99;
localparam signed [DEBIT:0]  W_8_x345 =  23'd125;
localparam signed [DEBIT:0]  W_8_x346 =  23'd84;
localparam signed [DEBIT:0]  W_8_x347 = - 23'd57;
localparam signed [DEBIT:0]  W_8_x348 = - 23'd3;
localparam signed [DEBIT:0]  W_8_x349 =  23'd402;
localparam signed [DEBIT:0]  W_8_x350 =  23'd495;
localparam signed [DEBIT:0]  W_8_x351 =  23'd155;
localparam signed [DEBIT:0]  W_8_x352 =  23'd82;
localparam signed [DEBIT:0]  W_8_x353 =  23'd38;
localparam signed [DEBIT:0]  W_8_x354 =  23'd44;
localparam signed [DEBIT:0]  W_8_x355 =  23'd49;
localparam signed [DEBIT:0]  W_8_x356 =  23'd221;
localparam signed [DEBIT:0]  W_8_x357 =  23'd26;
localparam signed [DEBIT:0]  W_8_x358 =  23'd97;
localparam signed [DEBIT:0]  W_8_x359 =  23'd24;
localparam signed [DEBIT:0]  W_8_x360 =  23'd237;
localparam signed [DEBIT:0]  W_8_x361 =  23'd583;
localparam signed [DEBIT:0]  W_8_x362 =  23'd850;
localparam signed [DEBIT:0]  W_8_x363 =  23'd917;
localparam signed [DEBIT:0]  W_8_x364 =  23'd934;
localparam signed [DEBIT:0]  W_8_x365 =  23'd938;
localparam signed [DEBIT:0]  W_8_x366 =  23'd941;
localparam signed [DEBIT:0]  W_8_x367 =  23'd883;
localparam signed [DEBIT:0]  W_8_x368 =  23'd705;
localparam signed [DEBIT:0]  W_8_x369 =  23'd437;
localparam signed [DEBIT:0]  W_8_x370 =  23'd71;
localparam signed [DEBIT:0]  W_8_x371 = - 23'd80;
localparam signed [DEBIT:0]  W_8_x372 = - 23'd84;
localparam signed [DEBIT:0]  W_8_x373 =  23'd17;
localparam signed [DEBIT:0]  W_8_x374 = - 23'd57;
localparam signed [DEBIT:0]  W_8_x375 = - 23'd139;
localparam signed [DEBIT:0]  W_8_x376 = - 23'd26;
localparam signed [DEBIT:0]  W_8_x377 =  23'd488;
localparam signed [DEBIT:0]  W_8_x378 =  23'd358;
localparam signed [DEBIT:0]  W_8_x379 = - 23'd38;
localparam signed [DEBIT:0]  W_8_x380 =  23'd114;
localparam signed [DEBIT:0]  W_8_x381 =  23'd141;
localparam signed [DEBIT:0]  W_8_x382 = - 23'd45;
localparam signed [DEBIT:0]  W_8_x383 = - 23'd98;
localparam signed [DEBIT:0]  W_8_x384 =  23'd11;
localparam signed [DEBIT:0]  W_8_x385 = - 23'd19;
localparam signed [DEBIT:0]  W_8_x386 = - 23'd25;
localparam signed [DEBIT:0]  W_8_x387 = - 23'd19;
localparam signed [DEBIT:0]  W_8_x388 =  23'd22;
localparam signed [DEBIT:0]  W_8_x389 =  23'd403;
localparam signed [DEBIT:0]  W_8_x390 =  23'd792;
localparam signed [DEBIT:0]  W_8_x391 =  23'd918;
localparam signed [DEBIT:0]  W_8_x392 =  23'd924;
localparam signed [DEBIT:0]  W_8_x393 =  23'd945;
localparam signed [DEBIT:0]  W_8_x394 =  23'd936;
localparam signed [DEBIT:0]  W_8_x395 =  23'd913;
localparam signed [DEBIT:0]  W_8_x396 =  23'd772;
localparam signed [DEBIT:0]  W_8_x397 =  23'd510;
localparam signed [DEBIT:0]  W_8_x398 =  23'd55;
localparam signed [DEBIT:0]  W_8_x399 = - 23'd310;
localparam signed [DEBIT:0]  W_8_x400 = - 23'd334;
localparam signed [DEBIT:0]  W_8_x401 = - 23'd310;
localparam signed [DEBIT:0]  W_8_x402 = - 23'd246;
localparam signed [DEBIT:0]  W_8_x403 = - 23'd163;
localparam signed [DEBIT:0]  W_8_x404 =  23'd190;
localparam signed [DEBIT:0]  W_8_x405 =  23'd364;
localparam signed [DEBIT:0]  W_8_x406 =  23'd191;
localparam signed [DEBIT:0]  W_8_x407 =  23'd40;
localparam signed [DEBIT:0]  W_8_x408 =  23'd97;
localparam signed [DEBIT:0]  W_8_x409 =  23'd85;
localparam signed [DEBIT:0]  W_8_x410 = - 23'd87;
localparam signed [DEBIT:0]  W_8_x411 = - 23'd198;
localparam signed [DEBIT:0]  W_8_x412 = - 23'd216;
localparam signed [DEBIT:0]  W_8_x413 = - 23'd157;
localparam signed [DEBIT:0]  W_8_x414 = - 23'd114;
localparam signed [DEBIT:0]  W_8_x415 = - 23'd100;
localparam signed [DEBIT:0]  W_8_x416 = - 23'd110;
localparam signed [DEBIT:0]  W_8_x417 =  23'd308;
localparam signed [DEBIT:0]  W_8_x418 =  23'd767;
localparam signed [DEBIT:0]  W_8_x419 =  23'd906;
localparam signed [DEBIT:0]  W_8_x420 =  23'd938;
localparam signed [DEBIT:0]  W_8_x421 =  23'd931;
localparam signed [DEBIT:0]  W_8_x422 =  23'd931;
localparam signed [DEBIT:0]  W_8_x423 =  23'd919;
localparam signed [DEBIT:0]  W_8_x424 =  23'd791;
localparam signed [DEBIT:0]  W_8_x425 =  23'd553;
localparam signed [DEBIT:0]  W_8_x426 = - 23'd6;
localparam signed [DEBIT:0]  W_8_x427 = - 23'd450;
localparam signed [DEBIT:0]  W_8_x428 = - 23'd501;
localparam signed [DEBIT:0]  W_8_x429 = - 23'd394;
localparam signed [DEBIT:0]  W_8_x430 = - 23'd266;
localparam signed [DEBIT:0]  W_8_x431 = - 23'd101;
localparam signed [DEBIT:0]  W_8_x432 =  23'd118;
localparam signed [DEBIT:0]  W_8_x433 =  23'd292;
localparam signed [DEBIT:0]  W_8_x434 =  23'd273;
localparam signed [DEBIT:0]  W_8_x435 =  23'd59;
localparam signed [DEBIT:0]  W_8_x436 =  23'd157;
localparam signed [DEBIT:0]  W_8_x437 =  23'd71;
localparam signed [DEBIT:0]  W_8_x438 = - 23'd224;
localparam signed [DEBIT:0]  W_8_x439 = - 23'd206;
localparam signed [DEBIT:0]  W_8_x440 = - 23'd259;
localparam signed [DEBIT:0]  W_8_x441 = - 23'd309;
localparam signed [DEBIT:0]  W_8_x442 = - 23'd176;
localparam signed [DEBIT:0]  W_8_x443 = - 23'd171;
localparam signed [DEBIT:0]  W_8_x444 = - 23'd145;
localparam signed [DEBIT:0]  W_8_x445 =  23'd239;
localparam signed [DEBIT:0]  W_8_x446 =  23'd722;
localparam signed [DEBIT:0]  W_8_x447 =  23'd881;
localparam signed [DEBIT:0]  W_8_x448 =  23'd938;
localparam signed [DEBIT:0]  W_8_x449 =  23'd940;
localparam signed [DEBIT:0]  W_8_x450 =  23'd938;
localparam signed [DEBIT:0]  W_8_x451 =  23'd900;
localparam signed [DEBIT:0]  W_8_x452 =  23'd789;
localparam signed [DEBIT:0]  W_8_x453 =  23'd509;
localparam signed [DEBIT:0]  W_8_x454 = - 23'd63;
localparam signed [DEBIT:0]  W_8_x455 = - 23'd440;
localparam signed [DEBIT:0]  W_8_x456 = - 23'd406;
localparam signed [DEBIT:0]  W_8_x457 = - 23'd133;
localparam signed [DEBIT:0]  W_8_x458 = - 23'd41;
localparam signed [DEBIT:0]  W_8_x459 =  23'd91;
localparam signed [DEBIT:0]  W_8_x460 =  23'd154;
localparam signed [DEBIT:0]  W_8_x461 =  23'd298;
localparam signed [DEBIT:0]  W_8_x462 =  23'd184;
localparam signed [DEBIT:0]  W_8_x463 = - 23'd28;
localparam signed [DEBIT:0]  W_8_x464 =  23'd178;
localparam signed [DEBIT:0]  W_8_x465 =  23'd100;
localparam signed [DEBIT:0]  W_8_x466 = - 23'd157;
localparam signed [DEBIT:0]  W_8_x467 = - 23'd375;
localparam signed [DEBIT:0]  W_8_x468 = - 23'd301;
localparam signed [DEBIT:0]  W_8_x469 = - 23'd203;
localparam signed [DEBIT:0]  W_8_x470 = - 23'd221;
localparam signed [DEBIT:0]  W_8_x471 = - 23'd186;
localparam signed [DEBIT:0]  W_8_x472 = - 23'd88;
localparam signed [DEBIT:0]  W_8_x473 =  23'd180;
localparam signed [DEBIT:0]  W_8_x474 =  23'd658;
localparam signed [DEBIT:0]  W_8_x475 =  23'd878;
localparam signed [DEBIT:0]  W_8_x476 =  23'd939;
localparam signed [DEBIT:0]  W_8_x477 =  23'd953;
localparam signed [DEBIT:0]  W_8_x478 =  23'd936;
localparam signed [DEBIT:0]  W_8_x479 =  23'd904;
localparam signed [DEBIT:0]  W_8_x480 =  23'd759;
localparam signed [DEBIT:0]  W_8_x481 =  23'd421;
localparam signed [DEBIT:0]  W_8_x482 = - 23'd101;
localparam signed [DEBIT:0]  W_8_x483 = - 23'd340;
localparam signed [DEBIT:0]  W_8_x484 = - 23'd159;
localparam signed [DEBIT:0]  W_8_x485 =  23'd220;
localparam signed [DEBIT:0]  W_8_x486 =  23'd311;
localparam signed [DEBIT:0]  W_8_x487 =  23'd271;
localparam signed [DEBIT:0]  W_8_x488 =  23'd333;
localparam signed [DEBIT:0]  W_8_x489 =  23'd449;
localparam signed [DEBIT:0]  W_8_x490 =  23'd104;
localparam signed [DEBIT:0]  W_8_x491 = - 23'd41;
localparam signed [DEBIT:0]  W_8_x492 = - 23'd103;
localparam signed [DEBIT:0]  W_8_x493 = - 23'd11;
localparam signed [DEBIT:0]  W_8_x494 = - 23'd61;
localparam signed [DEBIT:0]  W_8_x495 = - 23'd265;
localparam signed [DEBIT:0]  W_8_x496 = - 23'd205;
localparam signed [DEBIT:0]  W_8_x497 = - 23'd121;
localparam signed [DEBIT:0]  W_8_x498 = - 23'd212;
localparam signed [DEBIT:0]  W_8_x499 = - 23'd143;
localparam signed [DEBIT:0]  W_8_x500 = - 23'd65;
localparam signed [DEBIT:0]  W_8_x501 =  23'd199;
localparam signed [DEBIT:0]  W_8_x502 =  23'd655;
localparam signed [DEBIT:0]  W_8_x503 =  23'd882;
localparam signed [DEBIT:0]  W_8_x504 =  23'd943;
localparam signed [DEBIT:0]  W_8_x505 =  23'd936;
localparam signed [DEBIT:0]  W_8_x506 =  23'd936;
localparam signed [DEBIT:0]  W_8_x507 =  23'd900;
localparam signed [DEBIT:0]  W_8_x508 =  23'd670;
localparam signed [DEBIT:0]  W_8_x509 =  23'd286;
localparam signed [DEBIT:0]  W_8_x510 = - 23'd59;
localparam signed [DEBIT:0]  W_8_x511 = - 23'd138;
localparam signed [DEBIT:0]  W_8_x512 =  23'd43;
localparam signed [DEBIT:0]  W_8_x513 =  23'd344;
localparam signed [DEBIT:0]  W_8_x514 =  23'd382;
localparam signed [DEBIT:0]  W_8_x515 =  23'd271;
localparam signed [DEBIT:0]  W_8_x516 =  23'd431;
localparam signed [DEBIT:0]  W_8_x517 =  23'd307;
localparam signed [DEBIT:0]  W_8_x518 =  23'd36;
localparam signed [DEBIT:0]  W_8_x519 = - 23'd267;
localparam signed [DEBIT:0]  W_8_x520 = - 23'd270;
localparam signed [DEBIT:0]  W_8_x521 = - 23'd168;
localparam signed [DEBIT:0]  W_8_x522 = - 23'd257;
localparam signed [DEBIT:0]  W_8_x523 = - 23'd289;
localparam signed [DEBIT:0]  W_8_x524 = - 23'd104;
localparam signed [DEBIT:0]  W_8_x525 =  23'd40;
localparam signed [DEBIT:0]  W_8_x526 = - 23'd199;
localparam signed [DEBIT:0]  W_8_x527 = - 23'd238;
localparam signed [DEBIT:0]  W_8_x528 = - 23'd80;
localparam signed [DEBIT:0]  W_8_x529 =  23'd242;
localparam signed [DEBIT:0]  W_8_x530 =  23'd717;
localparam signed [DEBIT:0]  W_8_x531 =  23'd910;
localparam signed [DEBIT:0]  W_8_x532 =  23'd944;
localparam signed [DEBIT:0]  W_8_x533 =  23'd936;
localparam signed [DEBIT:0]  W_8_x534 =  23'd930;
localparam signed [DEBIT:0]  W_8_x535 =  23'd883;
localparam signed [DEBIT:0]  W_8_x536 =  23'd566;
localparam signed [DEBIT:0]  W_8_x537 =  23'd182;
localparam signed [DEBIT:0]  W_8_x538 =  23'd0;
localparam signed [DEBIT:0]  W_8_x539 = - 23'd90;
localparam signed [DEBIT:0]  W_8_x540 =  23'd38;
localparam signed [DEBIT:0]  W_8_x541 =  23'd195;
localparam signed [DEBIT:0]  W_8_x542 =  23'd182;
localparam signed [DEBIT:0]  W_8_x543 =  23'd85;
localparam signed [DEBIT:0]  W_8_x544 =  23'd33;
localparam signed [DEBIT:0]  W_8_x545 =  23'd36;
localparam signed [DEBIT:0]  W_8_x546 = - 23'd264;
localparam signed [DEBIT:0]  W_8_x547 = - 23'd372;
localparam signed [DEBIT:0]  W_8_x548 = - 23'd196;
localparam signed [DEBIT:0]  W_8_x549 = - 23'd192;
localparam signed [DEBIT:0]  W_8_x550 = - 23'd259;
localparam signed [DEBIT:0]  W_8_x551 = - 23'd315;
localparam signed [DEBIT:0]  W_8_x552 = - 23'd148;
localparam signed [DEBIT:0]  W_8_x553 = - 23'd36;
localparam signed [DEBIT:0]  W_8_x554 = - 23'd290;
localparam signed [DEBIT:0]  W_8_x555 = - 23'd292;
localparam signed [DEBIT:0]  W_8_x556 = - 23'd54;
localparam signed [DEBIT:0]  W_8_x557 =  23'd348;
localparam signed [DEBIT:0]  W_8_x558 =  23'd736;
localparam signed [DEBIT:0]  W_8_x559 =  23'd894;
localparam signed [DEBIT:0]  W_8_x560 =  23'd933;
localparam signed [DEBIT:0]  W_8_x561 =  23'd940;
localparam signed [DEBIT:0]  W_8_x562 =  23'd934;
localparam signed [DEBIT:0]  W_8_x563 =  23'd871;
localparam signed [DEBIT:0]  W_8_x564 =  23'd534;
localparam signed [DEBIT:0]  W_8_x565 =  23'd80;
localparam signed [DEBIT:0]  W_8_x566 = - 23'd22;
localparam signed [DEBIT:0]  W_8_x567 = - 23'd81;
localparam signed [DEBIT:0]  W_8_x568 =  23'd29;
localparam signed [DEBIT:0]  W_8_x569 =  23'd9;
localparam signed [DEBIT:0]  W_8_x570 =  23'd13;
localparam signed [DEBIT:0]  W_8_x571 = - 23'd44;
localparam signed [DEBIT:0]  W_8_x572 = - 23'd243;
localparam signed [DEBIT:0]  W_8_x573 = - 23'd156;
localparam signed [DEBIT:0]  W_8_x574 = - 23'd258;
localparam signed [DEBIT:0]  W_8_x575 = - 23'd295;
localparam signed [DEBIT:0]  W_8_x576 = - 23'd192;
localparam signed [DEBIT:0]  W_8_x577 = - 23'd316;
localparam signed [DEBIT:0]  W_8_x578 = - 23'd263;
localparam signed [DEBIT:0]  W_8_x579 = - 23'd271;
localparam signed [DEBIT:0]  W_8_x580 = - 23'd186;
localparam signed [DEBIT:0]  W_8_x581 = - 23'd201;
localparam signed [DEBIT:0]  W_8_x582 = - 23'd282;
localparam signed [DEBIT:0]  W_8_x583 = - 23'd270;
localparam signed [DEBIT:0]  W_8_x584 =  23'd28;
localparam signed [DEBIT:0]  W_8_x585 =  23'd387;
localparam signed [DEBIT:0]  W_8_x586 =  23'd759;
localparam signed [DEBIT:0]  W_8_x587 =  23'd887;
localparam signed [DEBIT:0]  W_8_x588 =  23'd938;
localparam signed [DEBIT:0]  W_8_x589 =  23'd929;
localparam signed [DEBIT:0]  W_8_x590 =  23'd933;
localparam signed [DEBIT:0]  W_8_x591 =  23'd855;
localparam signed [DEBIT:0]  W_8_x592 =  23'd593;
localparam signed [DEBIT:0]  W_8_x593 =  23'd115;
localparam signed [DEBIT:0]  W_8_x594 = - 23'd67;
localparam signed [DEBIT:0]  W_8_x595 = - 23'd145;
localparam signed [DEBIT:0]  W_8_x596 = - 23'd155;
localparam signed [DEBIT:0]  W_8_x597 = - 23'd69;
localparam signed [DEBIT:0]  W_8_x598 = - 23'd54;
localparam signed [DEBIT:0]  W_8_x599 = - 23'd94;
localparam signed [DEBIT:0]  W_8_x600 = - 23'd70;
localparam signed [DEBIT:0]  W_8_x601 = - 23'd18;
localparam signed [DEBIT:0]  W_8_x602 =  23'd33;
localparam signed [DEBIT:0]  W_8_x603 = - 23'd80;
localparam signed [DEBIT:0]  W_8_x604 = - 23'd38;
localparam signed [DEBIT:0]  W_8_x605 = - 23'd173;
localparam signed [DEBIT:0]  W_8_x606 = - 23'd122;
localparam signed [DEBIT:0]  W_8_x607 = - 23'd160;
localparam signed [DEBIT:0]  W_8_x608 = - 23'd183;
localparam signed [DEBIT:0]  W_8_x609 = - 23'd275;
localparam signed [DEBIT:0]  W_8_x610 = - 23'd339;
localparam signed [DEBIT:0]  W_8_x611 = - 23'd200;
localparam signed [DEBIT:0]  W_8_x612 =  23'd204;
localparam signed [DEBIT:0]  W_8_x613 =  23'd537;
localparam signed [DEBIT:0]  W_8_x614 =  23'd813;
localparam signed [DEBIT:0]  W_8_x615 =  23'd906;
localparam signed [DEBIT:0]  W_8_x616 =  23'd938;
localparam signed [DEBIT:0]  W_8_x617 =  23'd940;
localparam signed [DEBIT:0]  W_8_x618 =  23'd945;
localparam signed [DEBIT:0]  W_8_x619 =  23'd894;
localparam signed [DEBIT:0]  W_8_x620 =  23'd688;
localparam signed [DEBIT:0]  W_8_x621 =  23'd327;
localparam signed [DEBIT:0]  W_8_x622 =  23'd0;
localparam signed [DEBIT:0]  W_8_x623 = - 23'd157;
localparam signed [DEBIT:0]  W_8_x624 = - 23'd165;
localparam signed [DEBIT:0]  W_8_x625 = - 23'd32;
localparam signed [DEBIT:0]  W_8_x626 = - 23'd50;
localparam signed [DEBIT:0]  W_8_x627 =  23'd35;
localparam signed [DEBIT:0]  W_8_x628 =  23'd213;
localparam signed [DEBIT:0]  W_8_x629 =  23'd405;
localparam signed [DEBIT:0]  W_8_x630 =  23'd407;
localparam signed [DEBIT:0]  W_8_x631 =  23'd259;
localparam signed [DEBIT:0]  W_8_x632 =  23'd168;
localparam signed [DEBIT:0]  W_8_x633 =  23'd59;
localparam signed [DEBIT:0]  W_8_x634 =  23'd70;
localparam signed [DEBIT:0]  W_8_x635 = - 23'd8;
localparam signed [DEBIT:0]  W_8_x636 = - 23'd162;
localparam signed [DEBIT:0]  W_8_x637 = - 23'd252;
localparam signed [DEBIT:0]  W_8_x638 = - 23'd178;
localparam signed [DEBIT:0]  W_8_x639 =  23'd93;
localparam signed [DEBIT:0]  W_8_x640 =  23'd474;
localparam signed [DEBIT:0]  W_8_x641 =  23'd714;
localparam signed [DEBIT:0]  W_8_x642 =  23'd880;
localparam signed [DEBIT:0]  W_8_x643 =  23'd936;
localparam signed [DEBIT:0]  W_8_x644 =  23'd943;
localparam signed [DEBIT:0]  W_8_x645 =  23'd945;
localparam signed [DEBIT:0]  W_8_x646 =  23'd928;
localparam signed [DEBIT:0]  W_8_x647 =  23'd914;
localparam signed [DEBIT:0]  W_8_x648 =  23'd821;
localparam signed [DEBIT:0]  W_8_x649 =  23'd524;
localparam signed [DEBIT:0]  W_8_x650 =  23'd140;
localparam signed [DEBIT:0]  W_8_x651 = - 23'd213;
localparam signed [DEBIT:0]  W_8_x652 = - 23'd276;
localparam signed [DEBIT:0]  W_8_x653 = - 23'd65;
localparam signed [DEBIT:0]  W_8_x654 = - 23'd19;
localparam signed [DEBIT:0]  W_8_x655 =  23'd12;
localparam signed [DEBIT:0]  W_8_x656 =  23'd147;
localparam signed [DEBIT:0]  W_8_x657 =  23'd382;
localparam signed [DEBIT:0]  W_8_x658 =  23'd512;
localparam signed [DEBIT:0]  W_8_x659 =  23'd459;
localparam signed [DEBIT:0]  W_8_x660 =  23'd382;
localparam signed [DEBIT:0]  W_8_x661 =  23'd417;
localparam signed [DEBIT:0]  W_8_x662 =  23'd303;
localparam signed [DEBIT:0]  W_8_x663 =  23'd105;
localparam signed [DEBIT:0]  W_8_x664 =  23'd123;
localparam signed [DEBIT:0]  W_8_x665 =  23'd136;
localparam signed [DEBIT:0]  W_8_x666 =  23'd276;
localparam signed [DEBIT:0]  W_8_x667 =  23'd499;
localparam signed [DEBIT:0]  W_8_x668 =  23'd738;
localparam signed [DEBIT:0]  W_8_x669 =  23'd865;
localparam signed [DEBIT:0]  W_8_x670 =  23'd925;
localparam signed [DEBIT:0]  W_8_x671 =  23'd942;
localparam signed [DEBIT:0]  W_8_x672 =  23'd942;
localparam signed [DEBIT:0]  W_8_x673 =  23'd951;
localparam signed [DEBIT:0]  W_8_x674 =  23'd948;
localparam signed [DEBIT:0]  W_8_x675 =  23'd932;
localparam signed [DEBIT:0]  W_8_x676 =  23'd879;
localparam signed [DEBIT:0]  W_8_x677 =  23'd736;
localparam signed [DEBIT:0]  W_8_x678 =  23'd494;
localparam signed [DEBIT:0]  W_8_x679 =  23'd247;
localparam signed [DEBIT:0]  W_8_x680 =  23'd3;
localparam signed [DEBIT:0]  W_8_x681 =  23'd24;
localparam signed [DEBIT:0]  W_8_x682 =  23'd93;
localparam signed [DEBIT:0]  W_8_x683 =  23'd28;
localparam signed [DEBIT:0]  W_8_x684 = - 23'd15;
localparam signed [DEBIT:0]  W_8_x685 = - 23'd67;
localparam signed [DEBIT:0]  W_8_x686 =  23'd1;
localparam signed [DEBIT:0]  W_8_x687 =  23'd69;
localparam signed [DEBIT:0]  W_8_x688 =  23'd204;
localparam signed [DEBIT:0]  W_8_x689 =  23'd277;
localparam signed [DEBIT:0]  W_8_x690 =  23'd175;
localparam signed [DEBIT:0]  W_8_x691 =  23'd244;
localparam signed [DEBIT:0]  W_8_x692 =  23'd381;
localparam signed [DEBIT:0]  W_8_x693 =  23'd461;
localparam signed [DEBIT:0]  W_8_x694 =  23'd573;
localparam signed [DEBIT:0]  W_8_x695 =  23'd726;
localparam signed [DEBIT:0]  W_8_x696 =  23'd847;
localparam signed [DEBIT:0]  W_8_x697 =  23'd917;
localparam signed [DEBIT:0]  W_8_x698 =  23'd928;
localparam signed [DEBIT:0]  W_8_x699 =  23'd936;
localparam signed [DEBIT:0]  W_8_x700 =  23'd933;
localparam signed [DEBIT:0]  W_8_x701 =  23'd947;
localparam signed [DEBIT:0]  W_8_x702 =  23'd937;
localparam signed [DEBIT:0]  W_8_x703 =  23'd932;
localparam signed [DEBIT:0]  W_8_x704 =  23'd937;
localparam signed [DEBIT:0]  W_8_x705 =  23'd873;
localparam signed [DEBIT:0]  W_8_x706 =  23'd807;
localparam signed [DEBIT:0]  W_8_x707 =  23'd673;
localparam signed [DEBIT:0]  W_8_x708 =  23'd488;
localparam signed [DEBIT:0]  W_8_x709 =  23'd255;
localparam signed [DEBIT:0]  W_8_x710 =  23'd58;
localparam signed [DEBIT:0]  W_8_x711 = - 23'd76;
localparam signed [DEBIT:0]  W_8_x712 = - 23'd89;
localparam signed [DEBIT:0]  W_8_x713 = - 23'd119;
localparam signed [DEBIT:0]  W_8_x714 = - 23'd121;
localparam signed [DEBIT:0]  W_8_x715 =  23'd15;
localparam signed [DEBIT:0]  W_8_x716 =  23'd131;
localparam signed [DEBIT:0]  W_8_x717 =  23'd153;
localparam signed [DEBIT:0]  W_8_x718 =  23'd281;
localparam signed [DEBIT:0]  W_8_x719 =  23'd367;
localparam signed [DEBIT:0]  W_8_x720 =  23'd515;
localparam signed [DEBIT:0]  W_8_x721 =  23'd644;
localparam signed [DEBIT:0]  W_8_x722 =  23'd772;
localparam signed [DEBIT:0]  W_8_x723 =  23'd844;
localparam signed [DEBIT:0]  W_8_x724 =  23'd901;
localparam signed [DEBIT:0]  W_8_x725 =  23'd932;
localparam signed [DEBIT:0]  W_8_x726 =  23'd936;
localparam signed [DEBIT:0]  W_8_x727 =  23'd940;
localparam signed [DEBIT:0]  W_8_x728 =  23'd948;
localparam signed [DEBIT:0]  W_8_x729 =  23'd942;
localparam signed [DEBIT:0]  W_8_x730 =  23'd949;
localparam signed [DEBIT:0]  W_8_x731 =  23'd938;
localparam signed [DEBIT:0]  W_8_x732 =  23'd945;
localparam signed [DEBIT:0]  W_8_x733 =  23'd926;
localparam signed [DEBIT:0]  W_8_x734 =  23'd910;
localparam signed [DEBIT:0]  W_8_x735 =  23'd838;
localparam signed [DEBIT:0]  W_8_x736 =  23'd794;
localparam signed [DEBIT:0]  W_8_x737 =  23'd715;
localparam signed [DEBIT:0]  W_8_x738 =  23'd645;
localparam signed [DEBIT:0]  W_8_x739 =  23'd585;
localparam signed [DEBIT:0]  W_8_x740 =  23'd535;
localparam signed [DEBIT:0]  W_8_x741 =  23'd514;
localparam signed [DEBIT:0]  W_8_x742 =  23'd493;
localparam signed [DEBIT:0]  W_8_x743 =  23'd510;
localparam signed [DEBIT:0]  W_8_x744 =  23'd525;
localparam signed [DEBIT:0]  W_8_x745 =  23'd524;
localparam signed [DEBIT:0]  W_8_x746 =  23'd543;
localparam signed [DEBIT:0]  W_8_x747 =  23'd593;
localparam signed [DEBIT:0]  W_8_x748 =  23'd693;
localparam signed [DEBIT:0]  W_8_x749 =  23'd805;
localparam signed [DEBIT:0]  W_8_x750 =  23'd841;
localparam signed [DEBIT:0]  W_8_x751 =  23'd903;
localparam signed [DEBIT:0]  W_8_x752 =  23'd940;
localparam signed [DEBIT:0]  W_8_x753 =  23'd940;
localparam signed [DEBIT:0]  W_8_x754 =  23'd934;
localparam signed [DEBIT:0]  W_8_x755 =  23'd954;
localparam signed [DEBIT:0]  W_8_x756 =  23'd941;
localparam signed [DEBIT:0]  W_8_x757 =  23'd936;
localparam signed [DEBIT:0]  W_8_x758 =  23'd940;
localparam signed [DEBIT:0]  W_8_x759 =  23'd931;
localparam signed [DEBIT:0]  W_8_x760 =  23'd939;
localparam signed [DEBIT:0]  W_8_x761 =  23'd943;
localparam signed [DEBIT:0]  W_8_x762 =  23'd927;
localparam signed [DEBIT:0]  W_8_x763 =  23'd918;
localparam signed [DEBIT:0]  W_8_x764 =  23'd924;
localparam signed [DEBIT:0]  W_8_x765 =  23'd918;
localparam signed [DEBIT:0]  W_8_x766 =  23'd920;
localparam signed [DEBIT:0]  W_8_x767 =  23'd911;
localparam signed [DEBIT:0]  W_8_x768 =  23'd869;
localparam signed [DEBIT:0]  W_8_x769 =  23'd833;
localparam signed [DEBIT:0]  W_8_x770 =  23'd838;
localparam signed [DEBIT:0]  W_8_x771 =  23'd824;
localparam signed [DEBIT:0]  W_8_x772 =  23'd839;
localparam signed [DEBIT:0]  W_8_x773 =  23'd823;
localparam signed [DEBIT:0]  W_8_x774 =  23'd816;
localparam signed [DEBIT:0]  W_8_x775 =  23'd817;
localparam signed [DEBIT:0]  W_8_x776 =  23'd865;
localparam signed [DEBIT:0]  W_8_x777 =  23'd901;
localparam signed [DEBIT:0]  W_8_x778 =  23'd919;
localparam signed [DEBIT:0]  W_8_x779 =  23'd938;
localparam signed [DEBIT:0]  W_8_x780 =  23'd942;
localparam signed [DEBIT:0]  W_8_x781 =  23'd940;
localparam signed [DEBIT:0]  W_8_x782 =  23'd932;
localparam signed [DEBIT:0]  W_8_x783 =  23'd940;
localparam signed [DEBIT:0]  W_8_x784 =  23'd936;
localparam signed [DEBIT:0]  W_9_x1 =  23'd962;
localparam signed [DEBIT:0]  W_9_x2 =  23'd972;
localparam signed [DEBIT:0]  W_9_x3 =  23'd967;
localparam signed [DEBIT:0]  W_9_x4 =  23'd969;
localparam signed [DEBIT:0]  W_9_x5 =  23'd955;
localparam signed [DEBIT:0]  W_9_x6 =  23'd959;
localparam signed [DEBIT:0]  W_9_x7 =  23'd973;
localparam signed [DEBIT:0]  W_9_x8 =  23'd957;
localparam signed [DEBIT:0]  W_9_x9 =  23'd961;
localparam signed [DEBIT:0]  W_9_x10 =  23'd965;
localparam signed [DEBIT:0]  W_9_x11 =  23'd952;
localparam signed [DEBIT:0]  W_9_x12 =  23'd959;
localparam signed [DEBIT:0]  W_9_x13 =  23'd954;
localparam signed [DEBIT:0]  W_9_x14 =  23'd943;
localparam signed [DEBIT:0]  W_9_x15 =  23'd955;
localparam signed [DEBIT:0]  W_9_x16 =  23'd959;
localparam signed [DEBIT:0]  W_9_x17 =  23'd965;
localparam signed [DEBIT:0]  W_9_x18 =  23'd956;
localparam signed [DEBIT:0]  W_9_x19 =  23'd969;
localparam signed [DEBIT:0]  W_9_x20 =  23'd962;
localparam signed [DEBIT:0]  W_9_x21 =  23'd966;
localparam signed [DEBIT:0]  W_9_x22 =  23'd953;
localparam signed [DEBIT:0]  W_9_x23 =  23'd954;
localparam signed [DEBIT:0]  W_9_x24 =  23'd960;
localparam signed [DEBIT:0]  W_9_x25 =  23'd963;
localparam signed [DEBIT:0]  W_9_x26 =  23'd958;
localparam signed [DEBIT:0]  W_9_x27 =  23'd972;
localparam signed [DEBIT:0]  W_9_x28 =  23'd962;
localparam signed [DEBIT:0]  W_9_x29 =  23'd968;
localparam signed [DEBIT:0]  W_9_x30 =  23'd959;
localparam signed [DEBIT:0]  W_9_x31 =  23'd971;
localparam signed [DEBIT:0]  W_9_x32 =  23'd972;
localparam signed [DEBIT:0]  W_9_x33 =  23'd950;
localparam signed [DEBIT:0]  W_9_x34 =  23'd963;
localparam signed [DEBIT:0]  W_9_x35 =  23'd954;
localparam signed [DEBIT:0]  W_9_x36 =  23'd956;
localparam signed [DEBIT:0]  W_9_x37 =  23'd947;
localparam signed [DEBIT:0]  W_9_x38 =  23'd935;
localparam signed [DEBIT:0]  W_9_x39 =  23'd928;
localparam signed [DEBIT:0]  W_9_x40 =  23'd928;
localparam signed [DEBIT:0]  W_9_x41 =  23'd928;
localparam signed [DEBIT:0]  W_9_x42 =  23'd933;
localparam signed [DEBIT:0]  W_9_x43 =  23'd911;
localparam signed [DEBIT:0]  W_9_x44 =  23'd919;
localparam signed [DEBIT:0]  W_9_x45 =  23'd914;
localparam signed [DEBIT:0]  W_9_x46 =  23'd929;
localparam signed [DEBIT:0]  W_9_x47 =  23'd943;
localparam signed [DEBIT:0]  W_9_x48 =  23'd949;
localparam signed [DEBIT:0]  W_9_x49 =  23'd963;
localparam signed [DEBIT:0]  W_9_x50 =  23'd970;
localparam signed [DEBIT:0]  W_9_x51 =  23'd961;
localparam signed [DEBIT:0]  W_9_x52 =  23'd962;
localparam signed [DEBIT:0]  W_9_x53 =  23'd959;
localparam signed [DEBIT:0]  W_9_x54 =  23'd958;
localparam signed [DEBIT:0]  W_9_x55 =  23'd959;
localparam signed [DEBIT:0]  W_9_x56 =  23'd961;
localparam signed [DEBIT:0]  W_9_x57 =  23'd962;
localparam signed [DEBIT:0]  W_9_x58 =  23'd956;
localparam signed [DEBIT:0]  W_9_x59 =  23'd956;
localparam signed [DEBIT:0]  W_9_x60 =  23'd960;
localparam signed [DEBIT:0]  W_9_x61 =  23'd959;
localparam signed [DEBIT:0]  W_9_x62 =  23'd956;
localparam signed [DEBIT:0]  W_9_x63 =  23'd952;
localparam signed [DEBIT:0]  W_9_x64 =  23'd937;
localparam signed [DEBIT:0]  W_9_x65 =  23'd891;
localparam signed [DEBIT:0]  W_9_x66 =  23'd868;
localparam signed [DEBIT:0]  W_9_x67 =  23'd841;
localparam signed [DEBIT:0]  W_9_x68 =  23'd810;
localparam signed [DEBIT:0]  W_9_x69 =  23'd778;
localparam signed [DEBIT:0]  W_9_x70 =  23'd763;
localparam signed [DEBIT:0]  W_9_x71 =  23'd714;
localparam signed [DEBIT:0]  W_9_x72 =  23'd697;
localparam signed [DEBIT:0]  W_9_x73 =  23'd688;
localparam signed [DEBIT:0]  W_9_x74 =  23'd751;
localparam signed [DEBIT:0]  W_9_x75 =  23'd801;
localparam signed [DEBIT:0]  W_9_x76 =  23'd843;
localparam signed [DEBIT:0]  W_9_x77 =  23'd907;
localparam signed [DEBIT:0]  W_9_x78 =  23'd927;
localparam signed [DEBIT:0]  W_9_x79 =  23'd946;
localparam signed [DEBIT:0]  W_9_x80 =  23'd957;
localparam signed [DEBIT:0]  W_9_x81 =  23'd965;
localparam signed [DEBIT:0]  W_9_x82 =  23'd960;
localparam signed [DEBIT:0]  W_9_x83 =  23'd965;
localparam signed [DEBIT:0]  W_9_x84 =  23'd959;
localparam signed [DEBIT:0]  W_9_x85 =  23'd968;
localparam signed [DEBIT:0]  W_9_x86 =  23'd959;
localparam signed [DEBIT:0]  W_9_x87 =  23'd962;
localparam signed [DEBIT:0]  W_9_x88 =  23'd966;
localparam signed [DEBIT:0]  W_9_x89 =  23'd966;
localparam signed [DEBIT:0]  W_9_x90 =  23'd945;
localparam signed [DEBIT:0]  W_9_x91 =  23'd927;
localparam signed [DEBIT:0]  W_9_x92 =  23'd847;
localparam signed [DEBIT:0]  W_9_x93 =  23'd768;
localparam signed [DEBIT:0]  W_9_x94 =  23'd677;
localparam signed [DEBIT:0]  W_9_x95 =  23'd601;
localparam signed [DEBIT:0]  W_9_x96 =  23'd522;
localparam signed [DEBIT:0]  W_9_x97 =  23'd507;
localparam signed [DEBIT:0]  W_9_x98 =  23'd533;
localparam signed [DEBIT:0]  W_9_x99 =  23'd472;
localparam signed [DEBIT:0]  W_9_x100 =  23'd382;
localparam signed [DEBIT:0]  W_9_x101 =  23'd388;
localparam signed [DEBIT:0]  W_9_x102 =  23'd456;
localparam signed [DEBIT:0]  W_9_x103 =  23'd548;
localparam signed [DEBIT:0]  W_9_x104 =  23'd638;
localparam signed [DEBIT:0]  W_9_x105 =  23'd747;
localparam signed [DEBIT:0]  W_9_x106 =  23'd847;
localparam signed [DEBIT:0]  W_9_x107 =  23'd910;
localparam signed [DEBIT:0]  W_9_x108 =  23'd938;
localparam signed [DEBIT:0]  W_9_x109 =  23'd952;
localparam signed [DEBIT:0]  W_9_x110 =  23'd965;
localparam signed [DEBIT:0]  W_9_x111 =  23'd959;
localparam signed [DEBIT:0]  W_9_x112 =  23'd957;
localparam signed [DEBIT:0]  W_9_x113 =  23'd960;
localparam signed [DEBIT:0]  W_9_x114 =  23'd962;
localparam signed [DEBIT:0]  W_9_x115 =  23'd943;
localparam signed [DEBIT:0]  W_9_x116 =  23'd971;
localparam signed [DEBIT:0]  W_9_x117 =  23'd960;
localparam signed [DEBIT:0]  W_9_x118 =  23'd908;
localparam signed [DEBIT:0]  W_9_x119 =  23'd815;
localparam signed [DEBIT:0]  W_9_x120 =  23'd698;
localparam signed [DEBIT:0]  W_9_x121 =  23'd529;
localparam signed [DEBIT:0]  W_9_x122 =  23'd410;
localparam signed [DEBIT:0]  W_9_x123 =  23'd317;
localparam signed [DEBIT:0]  W_9_x124 =  23'd265;
localparam signed [DEBIT:0]  W_9_x125 =  23'd160;
localparam signed [DEBIT:0]  W_9_x126 =  23'd136;
localparam signed [DEBIT:0]  W_9_x127 =  23'd93;
localparam signed [DEBIT:0]  W_9_x128 = - 23'd12;
localparam signed [DEBIT:0]  W_9_x129 = - 23'd71;
localparam signed [DEBIT:0]  W_9_x130 =  23'd18;
localparam signed [DEBIT:0]  W_9_x131 =  23'd131;
localparam signed [DEBIT:0]  W_9_x132 =  23'd269;
localparam signed [DEBIT:0]  W_9_x133 =  23'd401;
localparam signed [DEBIT:0]  W_9_x134 =  23'd554;
localparam signed [DEBIT:0]  W_9_x135 =  23'd691;
localparam signed [DEBIT:0]  W_9_x136 =  23'd827;
localparam signed [DEBIT:0]  W_9_x137 =  23'd915;
localparam signed [DEBIT:0]  W_9_x138 =  23'd950;
localparam signed [DEBIT:0]  W_9_x139 =  23'd961;
localparam signed [DEBIT:0]  W_9_x140 =  23'd963;
localparam signed [DEBIT:0]  W_9_x141 =  23'd964;
localparam signed [DEBIT:0]  W_9_x142 =  23'd958;
localparam signed [DEBIT:0]  W_9_x143 =  23'd953;
localparam signed [DEBIT:0]  W_9_x144 =  23'd955;
localparam signed [DEBIT:0]  W_9_x145 =  23'd889;
localparam signed [DEBIT:0]  W_9_x146 =  23'd720;
localparam signed [DEBIT:0]  W_9_x147 =  23'd447;
localparam signed [DEBIT:0]  W_9_x148 =  23'd263;
localparam signed [DEBIT:0]  W_9_x149 =  23'd110;
localparam signed [DEBIT:0]  W_9_x150 = - 23'd10;
localparam signed [DEBIT:0]  W_9_x151 = - 23'd66;
localparam signed [DEBIT:0]  W_9_x152 = - 23'd30;
localparam signed [DEBIT:0]  W_9_x153 =  23'd17;
localparam signed [DEBIT:0]  W_9_x154 = - 23'd85;
localparam signed [DEBIT:0]  W_9_x155 = - 23'd191;
localparam signed [DEBIT:0]  W_9_x156 = - 23'd346;
localparam signed [DEBIT:0]  W_9_x157 = - 23'd418;
localparam signed [DEBIT:0]  W_9_x158 = - 23'd435;
localparam signed [DEBIT:0]  W_9_x159 = - 23'd437;
localparam signed [DEBIT:0]  W_9_x160 = - 23'd326;
localparam signed [DEBIT:0]  W_9_x161 = - 23'd196;
localparam signed [DEBIT:0]  W_9_x162 = - 23'd19;
localparam signed [DEBIT:0]  W_9_x163 =  23'd210;
localparam signed [DEBIT:0]  W_9_x164 =  23'd414;
localparam signed [DEBIT:0]  W_9_x165 =  23'd660;
localparam signed [DEBIT:0]  W_9_x166 =  23'd864;
localparam signed [DEBIT:0]  W_9_x167 =  23'd953;
localparam signed [DEBIT:0]  W_9_x168 =  23'd958;
localparam signed [DEBIT:0]  W_9_x169 =  23'd955;
localparam signed [DEBIT:0]  W_9_x170 =  23'd968;
localparam signed [DEBIT:0]  W_9_x171 =  23'd958;
localparam signed [DEBIT:0]  W_9_x172 =  23'd884;
localparam signed [DEBIT:0]  W_9_x173 =  23'd686;
localparam signed [DEBIT:0]  W_9_x174 =  23'd396;
localparam signed [DEBIT:0]  W_9_x175 =  23'd69;
localparam signed [DEBIT:0]  W_9_x176 = - 23'd241;
localparam signed [DEBIT:0]  W_9_x177 = - 23'd358;
localparam signed [DEBIT:0]  W_9_x178 = - 23'd358;
localparam signed [DEBIT:0]  W_9_x179 = - 23'd226;
localparam signed [DEBIT:0]  W_9_x180 =  23'd72;
localparam signed [DEBIT:0]  W_9_x181 =  23'd239;
localparam signed [DEBIT:0]  W_9_x182 =  23'd349;
localparam signed [DEBIT:0]  W_9_x183 =  23'd470;
localparam signed [DEBIT:0]  W_9_x184 =  23'd349;
localparam signed [DEBIT:0]  W_9_x185 =  23'd442;
localparam signed [DEBIT:0]  W_9_x186 =  23'd490;
localparam signed [DEBIT:0]  W_9_x187 =  23'd285;
localparam signed [DEBIT:0]  W_9_x188 = - 23'd16;
localparam signed [DEBIT:0]  W_9_x189 = - 23'd311;
localparam signed [DEBIT:0]  W_9_x190 = - 23'd422;
localparam signed [DEBIT:0]  W_9_x191 = - 23'd281;
localparam signed [DEBIT:0]  W_9_x192 = - 23'd26;
localparam signed [DEBIT:0]  W_9_x193 =  23'd296;
localparam signed [DEBIT:0]  W_9_x194 =  23'd663;
localparam signed [DEBIT:0]  W_9_x195 =  23'd904;
localparam signed [DEBIT:0]  W_9_x196 =  23'd952;
localparam signed [DEBIT:0]  W_9_x197 =  23'd964;
localparam signed [DEBIT:0]  W_9_x198 =  23'd945;
localparam signed [DEBIT:0]  W_9_x199 =  23'd921;
localparam signed [DEBIT:0]  W_9_x200 =  23'd746;
localparam signed [DEBIT:0]  W_9_x201 =  23'd425;
localparam signed [DEBIT:0]  W_9_x202 = - 23'd9;
localparam signed [DEBIT:0]  W_9_x203 = - 23'd351;
localparam signed [DEBIT:0]  W_9_x204 = - 23'd539;
localparam signed [DEBIT:0]  W_9_x205 = - 23'd327;
localparam signed [DEBIT:0]  W_9_x206 = - 23'd247;
localparam signed [DEBIT:0]  W_9_x207 = - 23'd46;
localparam signed [DEBIT:0]  W_9_x208 =  23'd75;
localparam signed [DEBIT:0]  W_9_x209 =  23'd260;
localparam signed [DEBIT:0]  W_9_x210 =  23'd392;
localparam signed [DEBIT:0]  W_9_x211 =  23'd589;
localparam signed [DEBIT:0]  W_9_x212 =  23'd697;
localparam signed [DEBIT:0]  W_9_x213 =  23'd595;
localparam signed [DEBIT:0]  W_9_x214 =  23'd321;
localparam signed [DEBIT:0]  W_9_x215 =  23'd156;
localparam signed [DEBIT:0]  W_9_x216 = - 23'd1;
localparam signed [DEBIT:0]  W_9_x217 = - 23'd226;
localparam signed [DEBIT:0]  W_9_x218 = - 23'd458;
localparam signed [DEBIT:0]  W_9_x219 = - 23'd531;
localparam signed [DEBIT:0]  W_9_x220 = - 23'd350;
localparam signed [DEBIT:0]  W_9_x221 =  23'd103;
localparam signed [DEBIT:0]  W_9_x222 =  23'd517;
localparam signed [DEBIT:0]  W_9_x223 =  23'd850;
localparam signed [DEBIT:0]  W_9_x224 =  23'd961;
localparam signed [DEBIT:0]  W_9_x225 =  23'd957;
localparam signed [DEBIT:0]  W_9_x226 =  23'd884;
localparam signed [DEBIT:0]  W_9_x227 =  23'd793;
localparam signed [DEBIT:0]  W_9_x228 =  23'd511;
localparam signed [DEBIT:0]  W_9_x229 =  23'd66;
localparam signed [DEBIT:0]  W_9_x230 = - 23'd377;
localparam signed [DEBIT:0]  W_9_x231 = - 23'd568;
localparam signed [DEBIT:0]  W_9_x232 = - 23'd500;
localparam signed [DEBIT:0]  W_9_x233 = - 23'd325;
localparam signed [DEBIT:0]  W_9_x234 = - 23'd192;
localparam signed [DEBIT:0]  W_9_x235 = - 23'd189;
localparam signed [DEBIT:0]  W_9_x236 = - 23'd179;
localparam signed [DEBIT:0]  W_9_x237 = - 23'd157;
localparam signed [DEBIT:0]  W_9_x238 =  23'd79;
localparam signed [DEBIT:0]  W_9_x239 =  23'd263;
localparam signed [DEBIT:0]  W_9_x240 =  23'd265;
localparam signed [DEBIT:0]  W_9_x241 =  23'd156;
localparam signed [DEBIT:0]  W_9_x242 = - 23'd113;
localparam signed [DEBIT:0]  W_9_x243 = - 23'd257;
localparam signed [DEBIT:0]  W_9_x244 = - 23'd250;
localparam signed [DEBIT:0]  W_9_x245 = - 23'd170;
localparam signed [DEBIT:0]  W_9_x246 = - 23'd400;
localparam signed [DEBIT:0]  W_9_x247 = - 23'd513;
localparam signed [DEBIT:0]  W_9_x248 = - 23'd324;
localparam signed [DEBIT:0]  W_9_x249 =  23'd149;
localparam signed [DEBIT:0]  W_9_x250 =  23'd529;
localparam signed [DEBIT:0]  W_9_x251 =  23'd850;
localparam signed [DEBIT:0]  W_9_x252 =  23'd954;
localparam signed [DEBIT:0]  W_9_x253 =  23'd957;
localparam signed [DEBIT:0]  W_9_x254 =  23'd874;
localparam signed [DEBIT:0]  W_9_x255 =  23'd723;
localparam signed [DEBIT:0]  W_9_x256 =  23'd399;
localparam signed [DEBIT:0]  W_9_x257 = - 23'd85;
localparam signed [DEBIT:0]  W_9_x258 = - 23'd492;
localparam signed [DEBIT:0]  W_9_x259 = - 23'd487;
localparam signed [DEBIT:0]  W_9_x260 = - 23'd301;
localparam signed [DEBIT:0]  W_9_x261 = - 23'd179;
localparam signed [DEBIT:0]  W_9_x262 = - 23'd152;
localparam signed [DEBIT:0]  W_9_x263 = - 23'd223;
localparam signed [DEBIT:0]  W_9_x264 = - 23'd83;
localparam signed [DEBIT:0]  W_9_x265 = - 23'd93;
localparam signed [DEBIT:0]  W_9_x266 = - 23'd97;
localparam signed [DEBIT:0]  W_9_x267 = - 23'd30;
localparam signed [DEBIT:0]  W_9_x268 =  23'd0;
localparam signed [DEBIT:0]  W_9_x269 = - 23'd214;
localparam signed [DEBIT:0]  W_9_x270 = - 23'd237;
localparam signed [DEBIT:0]  W_9_x271 = - 23'd217;
localparam signed [DEBIT:0]  W_9_x272 = - 23'd194;
localparam signed [DEBIT:0]  W_9_x273 = - 23'd113;
localparam signed [DEBIT:0]  W_9_x274 = - 23'd207;
localparam signed [DEBIT:0]  W_9_x275 = - 23'd333;
localparam signed [DEBIT:0]  W_9_x276 = - 23'd144;
localparam signed [DEBIT:0]  W_9_x277 =  23'd275;
localparam signed [DEBIT:0]  W_9_x278 =  23'd633;
localparam signed [DEBIT:0]  W_9_x279 =  23'd861;
localparam signed [DEBIT:0]  W_9_x280 =  23'd944;
localparam signed [DEBIT:0]  W_9_x281 =  23'd967;
localparam signed [DEBIT:0]  W_9_x282 =  23'd878;
localparam signed [DEBIT:0]  W_9_x283 =  23'd706;
localparam signed [DEBIT:0]  W_9_x284 =  23'd361;
localparam signed [DEBIT:0]  W_9_x285 = - 23'd88;
localparam signed [DEBIT:0]  W_9_x286 = - 23'd295;
localparam signed [DEBIT:0]  W_9_x287 = - 23'd263;
localparam signed [DEBIT:0]  W_9_x288 = - 23'd6;
localparam signed [DEBIT:0]  W_9_x289 =  23'd105;
localparam signed [DEBIT:0]  W_9_x290 = - 23'd46;
localparam signed [DEBIT:0]  W_9_x291 = - 23'd56;
localparam signed [DEBIT:0]  W_9_x292 =  23'd67;
localparam signed [DEBIT:0]  W_9_x293 = - 23'd59;
localparam signed [DEBIT:0]  W_9_x294 = - 23'd194;
localparam signed [DEBIT:0]  W_9_x295 = - 23'd273;
localparam signed [DEBIT:0]  W_9_x296 = - 23'd284;
localparam signed [DEBIT:0]  W_9_x297 = - 23'd273;
localparam signed [DEBIT:0]  W_9_x298 = - 23'd208;
localparam signed [DEBIT:0]  W_9_x299 = - 23'd150;
localparam signed [DEBIT:0]  W_9_x300 =  23'd24;
localparam signed [DEBIT:0]  W_9_x301 = - 23'd32;
localparam signed [DEBIT:0]  W_9_x302 = - 23'd47;
localparam signed [DEBIT:0]  W_9_x303 = - 23'd101;
localparam signed [DEBIT:0]  W_9_x304 =  23'd29;
localparam signed [DEBIT:0]  W_9_x305 =  23'd394;
localparam signed [DEBIT:0]  W_9_x306 =  23'd698;
localparam signed [DEBIT:0]  W_9_x307 =  23'd885;
localparam signed [DEBIT:0]  W_9_x308 =  23'd949;
localparam signed [DEBIT:0]  W_9_x309 =  23'd958;
localparam signed [DEBIT:0]  W_9_x310 =  23'd907;
localparam signed [DEBIT:0]  W_9_x311 =  23'd714;
localparam signed [DEBIT:0]  W_9_x312 =  23'd383;
localparam signed [DEBIT:0]  W_9_x313 =  23'd46;
localparam signed [DEBIT:0]  W_9_x314 = - 23'd67;
localparam signed [DEBIT:0]  W_9_x315 = - 23'd26;
localparam signed [DEBIT:0]  W_9_x316 =  23'd227;
localparam signed [DEBIT:0]  W_9_x317 =  23'd276;
localparam signed [DEBIT:0]  W_9_x318 =  23'd110;
localparam signed [DEBIT:0]  W_9_x319 =  23'd126;
localparam signed [DEBIT:0]  W_9_x320 =  23'd102;
localparam signed [DEBIT:0]  W_9_x321 = - 23'd71;
localparam signed [DEBIT:0]  W_9_x322 = - 23'd293;
localparam signed [DEBIT:0]  W_9_x323 = - 23'd257;
localparam signed [DEBIT:0]  W_9_x324 =  23'd64;
localparam signed [DEBIT:0]  W_9_x325 =  23'd73;
localparam signed [DEBIT:0]  W_9_x326 =  23'd134;
localparam signed [DEBIT:0]  W_9_x327 =  23'd20;
localparam signed [DEBIT:0]  W_9_x328 =  23'd182;
localparam signed [DEBIT:0]  W_9_x329 =  23'd240;
localparam signed [DEBIT:0]  W_9_x330 =  23'd119;
localparam signed [DEBIT:0]  W_9_x331 =  23'd2;
localparam signed [DEBIT:0]  W_9_x332 =  23'd165;
localparam signed [DEBIT:0]  W_9_x333 =  23'd519;
localparam signed [DEBIT:0]  W_9_x334 =  23'd781;
localparam signed [DEBIT:0]  W_9_x335 =  23'd891;
localparam signed [DEBIT:0]  W_9_x336 =  23'd957;
localparam signed [DEBIT:0]  W_9_x337 =  23'd964;
localparam signed [DEBIT:0]  W_9_x338 =  23'd920;
localparam signed [DEBIT:0]  W_9_x339 =  23'd770;
localparam signed [DEBIT:0]  W_9_x340 =  23'd526;
localparam signed [DEBIT:0]  W_9_x341 =  23'd285;
localparam signed [DEBIT:0]  W_9_x342 =  23'd173;
localparam signed [DEBIT:0]  W_9_x343 =  23'd227;
localparam signed [DEBIT:0]  W_9_x344 =  23'd291;
localparam signed [DEBIT:0]  W_9_x345 =  23'd230;
localparam signed [DEBIT:0]  W_9_x346 =  23'd211;
localparam signed [DEBIT:0]  W_9_x347 =  23'd226;
localparam signed [DEBIT:0]  W_9_x348 =  23'd123;
localparam signed [DEBIT:0]  W_9_x349 = - 23'd40;
localparam signed [DEBIT:0]  W_9_x350 = - 23'd120;
localparam signed [DEBIT:0]  W_9_x351 =  23'd28;
localparam signed [DEBIT:0]  W_9_x352 =  23'd234;
localparam signed [DEBIT:0]  W_9_x353 =  23'd182;
localparam signed [DEBIT:0]  W_9_x354 =  23'd225;
localparam signed [DEBIT:0]  W_9_x355 =  23'd166;
localparam signed [DEBIT:0]  W_9_x356 =  23'd305;
localparam signed [DEBIT:0]  W_9_x357 =  23'd193;
localparam signed [DEBIT:0]  W_9_x358 =  23'd136;
localparam signed [DEBIT:0]  W_9_x359 =  23'd69;
localparam signed [DEBIT:0]  W_9_x360 =  23'd211;
localparam signed [DEBIT:0]  W_9_x361 =  23'd482;
localparam signed [DEBIT:0]  W_9_x362 =  23'd791;
localparam signed [DEBIT:0]  W_9_x363 =  23'd898;
localparam signed [DEBIT:0]  W_9_x364 =  23'd948;
localparam signed [DEBIT:0]  W_9_x365 =  23'd964;
localparam signed [DEBIT:0]  W_9_x366 =  23'd944;
localparam signed [DEBIT:0]  W_9_x367 =  23'd858;
localparam signed [DEBIT:0]  W_9_x368 =  23'd700;
localparam signed [DEBIT:0]  W_9_x369 =  23'd503;
localparam signed [DEBIT:0]  W_9_x370 =  23'd389;
localparam signed [DEBIT:0]  W_9_x371 =  23'd339;
localparam signed [DEBIT:0]  W_9_x372 =  23'd308;
localparam signed [DEBIT:0]  W_9_x373 =  23'd208;
localparam signed [DEBIT:0]  W_9_x374 =  23'd228;
localparam signed [DEBIT:0]  W_9_x375 =  23'd257;
localparam signed [DEBIT:0]  W_9_x376 =  23'd110;
localparam signed [DEBIT:0]  W_9_x377 =  23'd32;
localparam signed [DEBIT:0]  W_9_x378 =  23'd78;
localparam signed [DEBIT:0]  W_9_x379 =  23'd114;
localparam signed [DEBIT:0]  W_9_x380 =  23'd228;
localparam signed [DEBIT:0]  W_9_x381 =  23'd199;
localparam signed [DEBIT:0]  W_9_x382 =  23'd160;
localparam signed [DEBIT:0]  W_9_x383 =  23'd219;
localparam signed [DEBIT:0]  W_9_x384 =  23'd260;
localparam signed [DEBIT:0]  W_9_x385 =  23'd85;
localparam signed [DEBIT:0]  W_9_x386 =  23'd37;
localparam signed [DEBIT:0]  W_9_x387 = - 23'd5;
localparam signed [DEBIT:0]  W_9_x388 =  23'd60;
localparam signed [DEBIT:0]  W_9_x389 =  23'd408;
localparam signed [DEBIT:0]  W_9_x390 =  23'd785;
localparam signed [DEBIT:0]  W_9_x391 =  23'd914;
localparam signed [DEBIT:0]  W_9_x392 =  23'd957;
localparam signed [DEBIT:0]  W_9_x393 =  23'd965;
localparam signed [DEBIT:0]  W_9_x394 =  23'd952;
localparam signed [DEBIT:0]  W_9_x395 =  23'd926;
localparam signed [DEBIT:0]  W_9_x396 =  23'd789;
localparam signed [DEBIT:0]  W_9_x397 =  23'd597;
localparam signed [DEBIT:0]  W_9_x398 =  23'd308;
localparam signed [DEBIT:0]  W_9_x399 =  23'd237;
localparam signed [DEBIT:0]  W_9_x400 =  23'd222;
localparam signed [DEBIT:0]  W_9_x401 =  23'd97;
localparam signed [DEBIT:0]  W_9_x402 =  23'd36;
localparam signed [DEBIT:0]  W_9_x403 =  23'd51;
localparam signed [DEBIT:0]  W_9_x404 =  23'd7;
localparam signed [DEBIT:0]  W_9_x405 =  23'd31;
localparam signed [DEBIT:0]  W_9_x406 =  23'd23;
localparam signed [DEBIT:0]  W_9_x407 =  23'd106;
localparam signed [DEBIT:0]  W_9_x408 =  23'd125;
localparam signed [DEBIT:0]  W_9_x409 =  23'd66;
localparam signed [DEBIT:0]  W_9_x410 =  23'd11;
localparam signed [DEBIT:0]  W_9_x411 =  23'd74;
localparam signed [DEBIT:0]  W_9_x412 =  23'd45;
localparam signed [DEBIT:0]  W_9_x413 = - 23'd28;
localparam signed [DEBIT:0]  W_9_x414 = - 23'd174;
localparam signed [DEBIT:0]  W_9_x415 = - 23'd123;
localparam signed [DEBIT:0]  W_9_x416 = - 23'd21;
localparam signed [DEBIT:0]  W_9_x417 =  23'd351;
localparam signed [DEBIT:0]  W_9_x418 =  23'd799;
localparam signed [DEBIT:0]  W_9_x419 =  23'd942;
localparam signed [DEBIT:0]  W_9_x420 =  23'd967;
localparam signed [DEBIT:0]  W_9_x421 =  23'd962;
localparam signed [DEBIT:0]  W_9_x422 =  23'd962;
localparam signed [DEBIT:0]  W_9_x423 =  23'd955;
localparam signed [DEBIT:0]  W_9_x424 =  23'd782;
localparam signed [DEBIT:0]  W_9_x425 =  23'd612;
localparam signed [DEBIT:0]  W_9_x426 =  23'd126;
localparam signed [DEBIT:0]  W_9_x427 = - 23'd73;
localparam signed [DEBIT:0]  W_9_x428 = - 23'd21;
localparam signed [DEBIT:0]  W_9_x429 =  23'd102;
localparam signed [DEBIT:0]  W_9_x430 =  23'd96;
localparam signed [DEBIT:0]  W_9_x431 =  23'd55;
localparam signed [DEBIT:0]  W_9_x432 =  23'd91;
localparam signed [DEBIT:0]  W_9_x433 =  23'd101;
localparam signed [DEBIT:0]  W_9_x434 = - 23'd123;
localparam signed [DEBIT:0]  W_9_x435 = - 23'd173;
localparam signed [DEBIT:0]  W_9_x436 = - 23'd64;
localparam signed [DEBIT:0]  W_9_x437 =  23'd58;
localparam signed [DEBIT:0]  W_9_x438 =  23'd102;
localparam signed [DEBIT:0]  W_9_x439 =  23'd7;
localparam signed [DEBIT:0]  W_9_x440 = - 23'd128;
localparam signed [DEBIT:0]  W_9_x441 = - 23'd173;
localparam signed [DEBIT:0]  W_9_x442 = - 23'd232;
localparam signed [DEBIT:0]  W_9_x443 = - 23'd193;
localparam signed [DEBIT:0]  W_9_x444 = - 23'd45;
localparam signed [DEBIT:0]  W_9_x445 =  23'd337;
localparam signed [DEBIT:0]  W_9_x446 =  23'd756;
localparam signed [DEBIT:0]  W_9_x447 =  23'd917;
localparam signed [DEBIT:0]  W_9_x448 =  23'd954;
localparam signed [DEBIT:0]  W_9_x449 =  23'd967;
localparam signed [DEBIT:0]  W_9_x450 =  23'd961;
localparam signed [DEBIT:0]  W_9_x451 =  23'd942;
localparam signed [DEBIT:0]  W_9_x452 =  23'd801;
localparam signed [DEBIT:0]  W_9_x453 =  23'd573;
localparam signed [DEBIT:0]  W_9_x454 =  23'd36;
localparam signed [DEBIT:0]  W_9_x455 = - 23'd201;
localparam signed [DEBIT:0]  W_9_x456 = - 23'd64;
localparam signed [DEBIT:0]  W_9_x457 =  23'd90;
localparam signed [DEBIT:0]  W_9_x458 =  23'd124;
localparam signed [DEBIT:0]  W_9_x459 =  23'd166;
localparam signed [DEBIT:0]  W_9_x460 =  23'd195;
localparam signed [DEBIT:0]  W_9_x461 =  23'd84;
localparam signed [DEBIT:0]  W_9_x462 = - 23'd137;
localparam signed [DEBIT:0]  W_9_x463 = - 23'd216;
localparam signed [DEBIT:0]  W_9_x464 =  23'd14;
localparam signed [DEBIT:0]  W_9_x465 =  23'd91;
localparam signed [DEBIT:0]  W_9_x466 =  23'd91;
localparam signed [DEBIT:0]  W_9_x467 = - 23'd127;
localparam signed [DEBIT:0]  W_9_x468 = - 23'd295;
localparam signed [DEBIT:0]  W_9_x469 = - 23'd256;
localparam signed [DEBIT:0]  W_9_x470 = - 23'd331;
localparam signed [DEBIT:0]  W_9_x471 = - 23'd176;
localparam signed [DEBIT:0]  W_9_x472 = - 23'd45;
localparam signed [DEBIT:0]  W_9_x473 =  23'd263;
localparam signed [DEBIT:0]  W_9_x474 =  23'd706;
localparam signed [DEBIT:0]  W_9_x475 =  23'd908;
localparam signed [DEBIT:0]  W_9_x476 =  23'd946;
localparam signed [DEBIT:0]  W_9_x477 =  23'd959;
localparam signed [DEBIT:0]  W_9_x478 =  23'd957;
localparam signed [DEBIT:0]  W_9_x479 =  23'd934;
localparam signed [DEBIT:0]  W_9_x480 =  23'd803;
localparam signed [DEBIT:0]  W_9_x481 =  23'd516;
localparam signed [DEBIT:0]  W_9_x482 =  23'd47;
localparam signed [DEBIT:0]  W_9_x483 = - 23'd115;
localparam signed [DEBIT:0]  W_9_x484 = - 23'd11;
localparam signed [DEBIT:0]  W_9_x485 =  23'd95;
localparam signed [DEBIT:0]  W_9_x486 =  23'd175;
localparam signed [DEBIT:0]  W_9_x487 =  23'd171;
localparam signed [DEBIT:0]  W_9_x488 =  23'd115;
localparam signed [DEBIT:0]  W_9_x489 =  23'd26;
localparam signed [DEBIT:0]  W_9_x490 = - 23'd104;
localparam signed [DEBIT:0]  W_9_x491 = - 23'd158;
localparam signed [DEBIT:0]  W_9_x492 =  23'd72;
localparam signed [DEBIT:0]  W_9_x493 =  23'd15;
localparam signed [DEBIT:0]  W_9_x494 = - 23'd48;
localparam signed [DEBIT:0]  W_9_x495 = - 23'd179;
localparam signed [DEBIT:0]  W_9_x496 = - 23'd246;
localparam signed [DEBIT:0]  W_9_x497 = - 23'd373;
localparam signed [DEBIT:0]  W_9_x498 = - 23'd435;
localparam signed [DEBIT:0]  W_9_x499 = - 23'd271;
localparam signed [DEBIT:0]  W_9_x500 = - 23'd76;
localparam signed [DEBIT:0]  W_9_x501 =  23'd265;
localparam signed [DEBIT:0]  W_9_x502 =  23'd750;
localparam signed [DEBIT:0]  W_9_x503 =  23'd921;
localparam signed [DEBIT:0]  W_9_x504 =  23'd962;
localparam signed [DEBIT:0]  W_9_x505 =  23'd967;
localparam signed [DEBIT:0]  W_9_x506 =  23'd958;
localparam signed [DEBIT:0]  W_9_x507 =  23'd924;
localparam signed [DEBIT:0]  W_9_x508 =  23'd747;
localparam signed [DEBIT:0]  W_9_x509 =  23'd470;
localparam signed [DEBIT:0]  W_9_x510 =  23'd38;
localparam signed [DEBIT:0]  W_9_x511 = - 23'd86;
localparam signed [DEBIT:0]  W_9_x512 = - 23'd101;
localparam signed [DEBIT:0]  W_9_x513 = - 23'd2;
localparam signed [DEBIT:0]  W_9_x514 = - 23'd5;
localparam signed [DEBIT:0]  W_9_x515 =  23'd18;
localparam signed [DEBIT:0]  W_9_x516 =  23'd36;
localparam signed [DEBIT:0]  W_9_x517 = - 23'd42;
localparam signed [DEBIT:0]  W_9_x518 = - 23'd129;
localparam signed [DEBIT:0]  W_9_x519 = - 23'd135;
localparam signed [DEBIT:0]  W_9_x520 = - 23'd167;
localparam signed [DEBIT:0]  W_9_x521 = - 23'd134;
localparam signed [DEBIT:0]  W_9_x522 = - 23'd260;
localparam signed [DEBIT:0]  W_9_x523 = - 23'd290;
localparam signed [DEBIT:0]  W_9_x524 = - 23'd185;
localparam signed [DEBIT:0]  W_9_x525 = - 23'd265;
localparam signed [DEBIT:0]  W_9_x526 = - 23'd481;
localparam signed [DEBIT:0]  W_9_x527 = - 23'd373;
localparam signed [DEBIT:0]  W_9_x528 = - 23'd83;
localparam signed [DEBIT:0]  W_9_x529 =  23'd383;
localparam signed [DEBIT:0]  W_9_x530 =  23'd814;
localparam signed [DEBIT:0]  W_9_x531 =  23'd933;
localparam signed [DEBIT:0]  W_9_x532 =  23'd961;
localparam signed [DEBIT:0]  W_9_x533 =  23'd967;
localparam signed [DEBIT:0]  W_9_x534 =  23'd954;
localparam signed [DEBIT:0]  W_9_x535 =  23'd884;
localparam signed [DEBIT:0]  W_9_x536 =  23'd672;
localparam signed [DEBIT:0]  W_9_x537 =  23'd408;
localparam signed [DEBIT:0]  W_9_x538 =  23'd55;
localparam signed [DEBIT:0]  W_9_x539 = - 23'd224;
localparam signed [DEBIT:0]  W_9_x540 = - 23'd295;
localparam signed [DEBIT:0]  W_9_x541 = - 23'd295;
localparam signed [DEBIT:0]  W_9_x542 = - 23'd319;
localparam signed [DEBIT:0]  W_9_x543 = - 23'd369;
localparam signed [DEBIT:0]  W_9_x544 = - 23'd286;
localparam signed [DEBIT:0]  W_9_x545 = - 23'd336;
localparam signed [DEBIT:0]  W_9_x546 = - 23'd254;
localparam signed [DEBIT:0]  W_9_x547 = - 23'd267;
localparam signed [DEBIT:0]  W_9_x548 = - 23'd346;
localparam signed [DEBIT:0]  W_9_x549 = - 23'd325;
localparam signed [DEBIT:0]  W_9_x550 = - 23'd349;
localparam signed [DEBIT:0]  W_9_x551 = - 23'd400;
localparam signed [DEBIT:0]  W_9_x552 = - 23'd215;
localparam signed [DEBIT:0]  W_9_x553 = - 23'd289;
localparam signed [DEBIT:0]  W_9_x554 = - 23'd576;
localparam signed [DEBIT:0]  W_9_x555 = - 23'd390;
localparam signed [DEBIT:0]  W_9_x556 =  23'd30;
localparam signed [DEBIT:0]  W_9_x557 =  23'd556;
localparam signed [DEBIT:0]  W_9_x558 =  23'd833;
localparam signed [DEBIT:0]  W_9_x559 =  23'd933;
localparam signed [DEBIT:0]  W_9_x560 =  23'd967;
localparam signed [DEBIT:0]  W_9_x561 =  23'd966;
localparam signed [DEBIT:0]  W_9_x562 =  23'd952;
localparam signed [DEBIT:0]  W_9_x563 =  23'd867;
localparam signed [DEBIT:0]  W_9_x564 =  23'd652;
localparam signed [DEBIT:0]  W_9_x565 =  23'd340;
localparam signed [DEBIT:0]  W_9_x566 =  23'd107;
localparam signed [DEBIT:0]  W_9_x567 = - 23'd220;
localparam signed [DEBIT:0]  W_9_x568 = - 23'd383;
localparam signed [DEBIT:0]  W_9_x569 = - 23'd433;
localparam signed [DEBIT:0]  W_9_x570 = - 23'd465;
localparam signed [DEBIT:0]  W_9_x571 = - 23'd464;
localparam signed [DEBIT:0]  W_9_x572 = - 23'd440;
localparam signed [DEBIT:0]  W_9_x573 = - 23'd505;
localparam signed [DEBIT:0]  W_9_x574 = - 23'd398;
localparam signed [DEBIT:0]  W_9_x575 = - 23'd377;
localparam signed [DEBIT:0]  W_9_x576 = - 23'd418;
localparam signed [DEBIT:0]  W_9_x577 = - 23'd285;
localparam signed [DEBIT:0]  W_9_x578 = - 23'd345;
localparam signed [DEBIT:0]  W_9_x579 = - 23'd349;
localparam signed [DEBIT:0]  W_9_x580 = - 23'd195;
localparam signed [DEBIT:0]  W_9_x581 = - 23'd425;
localparam signed [DEBIT:0]  W_9_x582 = - 23'd525;
localparam signed [DEBIT:0]  W_9_x583 = - 23'd262;
localparam signed [DEBIT:0]  W_9_x584 =  23'd174;
localparam signed [DEBIT:0]  W_9_x585 =  23'd655;
localparam signed [DEBIT:0]  W_9_x586 =  23'd871;
localparam signed [DEBIT:0]  W_9_x587 =  23'd941;
localparam signed [DEBIT:0]  W_9_x588 =  23'd961;
localparam signed [DEBIT:0]  W_9_x589 =  23'd959;
localparam signed [DEBIT:0]  W_9_x590 =  23'd962;
localparam signed [DEBIT:0]  W_9_x591 =  23'd885;
localparam signed [DEBIT:0]  W_9_x592 =  23'd676;
localparam signed [DEBIT:0]  W_9_x593 =  23'd412;
localparam signed [DEBIT:0]  W_9_x594 =  23'd115;
localparam signed [DEBIT:0]  W_9_x595 = - 23'd213;
localparam signed [DEBIT:0]  W_9_x596 = - 23'd395;
localparam signed [DEBIT:0]  W_9_x597 = - 23'd333;
localparam signed [DEBIT:0]  W_9_x598 = - 23'd255;
localparam signed [DEBIT:0]  W_9_x599 = - 23'd186;
localparam signed [DEBIT:0]  W_9_x600 = - 23'd278;
localparam signed [DEBIT:0]  W_9_x601 = - 23'd259;
localparam signed [DEBIT:0]  W_9_x602 = - 23'd261;
localparam signed [DEBIT:0]  W_9_x603 = - 23'd137;
localparam signed [DEBIT:0]  W_9_x604 = - 23'd146;
localparam signed [DEBIT:0]  W_9_x605 = - 23'd243;
localparam signed [DEBIT:0]  W_9_x606 = - 23'd260;
localparam signed [DEBIT:0]  W_9_x607 = - 23'd221;
localparam signed [DEBIT:0]  W_9_x608 = - 23'd230;
localparam signed [DEBIT:0]  W_9_x609 = - 23'd363;
localparam signed [DEBIT:0]  W_9_x610 = - 23'd399;
localparam signed [DEBIT:0]  W_9_x611 = - 23'd98;
localparam signed [DEBIT:0]  W_9_x612 =  23'd425;
localparam signed [DEBIT:0]  W_9_x613 =  23'd725;
localparam signed [DEBIT:0]  W_9_x614 =  23'd881;
localparam signed [DEBIT:0]  W_9_x615 =  23'd939;
localparam signed [DEBIT:0]  W_9_x616 =  23'd968;
localparam signed [DEBIT:0]  W_9_x617 =  23'd963;
localparam signed [DEBIT:0]  W_9_x618 =  23'd961;
localparam signed [DEBIT:0]  W_9_x619 =  23'd908;
localparam signed [DEBIT:0]  W_9_x620 =  23'd773;
localparam signed [DEBIT:0]  W_9_x621 =  23'd516;
localparam signed [DEBIT:0]  W_9_x622 =  23'd214;
localparam signed [DEBIT:0]  W_9_x623 = - 23'd131;
localparam signed [DEBIT:0]  W_9_x624 = - 23'd369;
localparam signed [DEBIT:0]  W_9_x625 = - 23'd232;
localparam signed [DEBIT:0]  W_9_x626 = - 23'd117;
localparam signed [DEBIT:0]  W_9_x627 = - 23'd5;
localparam signed [DEBIT:0]  W_9_x628 = - 23'd26;
localparam signed [DEBIT:0]  W_9_x629 =  23'd9;
localparam signed [DEBIT:0]  W_9_x630 = - 23'd24;
localparam signed [DEBIT:0]  W_9_x631 = - 23'd22;
localparam signed [DEBIT:0]  W_9_x632 = - 23'd130;
localparam signed [DEBIT:0]  W_9_x633 = - 23'd141;
localparam signed [DEBIT:0]  W_9_x634 = - 23'd199;
localparam signed [DEBIT:0]  W_9_x635 = - 23'd241;
localparam signed [DEBIT:0]  W_9_x636 = - 23'd277;
localparam signed [DEBIT:0]  W_9_x637 = - 23'd175;
localparam signed [DEBIT:0]  W_9_x638 = - 23'd101;
localparam signed [DEBIT:0]  W_9_x639 =  23'd223;
localparam signed [DEBIT:0]  W_9_x640 =  23'd663;
localparam signed [DEBIT:0]  W_9_x641 =  23'd872;
localparam signed [DEBIT:0]  W_9_x642 =  23'd931;
localparam signed [DEBIT:0]  W_9_x643 =  23'd960;
localparam signed [DEBIT:0]  W_9_x644 =  23'd966;
localparam signed [DEBIT:0]  W_9_x645 =  23'd961;
localparam signed [DEBIT:0]  W_9_x646 =  23'd966;
localparam signed [DEBIT:0]  W_9_x647 =  23'd943;
localparam signed [DEBIT:0]  W_9_x648 =  23'd880;
localparam signed [DEBIT:0]  W_9_x649 =  23'd691;
localparam signed [DEBIT:0]  W_9_x650 =  23'd451;
localparam signed [DEBIT:0]  W_9_x651 =  23'd56;
localparam signed [DEBIT:0]  W_9_x652 = - 23'd136;
localparam signed [DEBIT:0]  W_9_x653 = - 23'd121;
localparam signed [DEBIT:0]  W_9_x654 = - 23'd260;
localparam signed [DEBIT:0]  W_9_x655 = - 23'd226;
localparam signed [DEBIT:0]  W_9_x656 = - 23'd137;
localparam signed [DEBIT:0]  W_9_x657 = - 23'd144;
localparam signed [DEBIT:0]  W_9_x658 = - 23'd197;
localparam signed [DEBIT:0]  W_9_x659 = - 23'd208;
localparam signed [DEBIT:0]  W_9_x660 = - 23'd141;
localparam signed [DEBIT:0]  W_9_x661 = - 23'd69;
localparam signed [DEBIT:0]  W_9_x662 = - 23'd106;
localparam signed [DEBIT:0]  W_9_x663 = - 23'd157;
localparam signed [DEBIT:0]  W_9_x664 =  23'd112;
localparam signed [DEBIT:0]  W_9_x665 =  23'd272;
localparam signed [DEBIT:0]  W_9_x666 =  23'd411;
localparam signed [DEBIT:0]  W_9_x667 =  23'd640;
localparam signed [DEBIT:0]  W_9_x668 =  23'd843;
localparam signed [DEBIT:0]  W_9_x669 =  23'd967;
localparam signed [DEBIT:0]  W_9_x670 =  23'd964;
localparam signed [DEBIT:0]  W_9_x671 =  23'd965;
localparam signed [DEBIT:0]  W_9_x672 =  23'd956;
localparam signed [DEBIT:0]  W_9_x673 =  23'd970;
localparam signed [DEBIT:0]  W_9_x674 =  23'd970;
localparam signed [DEBIT:0]  W_9_x675 =  23'd946;
localparam signed [DEBIT:0]  W_9_x676 =  23'd926;
localparam signed [DEBIT:0]  W_9_x677 =  23'd827;
localparam signed [DEBIT:0]  W_9_x678 =  23'd679;
localparam signed [DEBIT:0]  W_9_x679 =  23'd451;
localparam signed [DEBIT:0]  W_9_x680 =  23'd284;
localparam signed [DEBIT:0]  W_9_x681 =  23'd161;
localparam signed [DEBIT:0]  W_9_x682 = - 23'd14;
localparam signed [DEBIT:0]  W_9_x683 = - 23'd57;
localparam signed [DEBIT:0]  W_9_x684 = - 23'd46;
localparam signed [DEBIT:0]  W_9_x685 = - 23'd100;
localparam signed [DEBIT:0]  W_9_x686 = - 23'd58;
localparam signed [DEBIT:0]  W_9_x687 = - 23'd35;
localparam signed [DEBIT:0]  W_9_x688 =  23'd75;
localparam signed [DEBIT:0]  W_9_x689 =  23'd94;
localparam signed [DEBIT:0]  W_9_x690 =  23'd256;
localparam signed [DEBIT:0]  W_9_x691 =  23'd365;
localparam signed [DEBIT:0]  W_9_x692 =  23'd635;
localparam signed [DEBIT:0]  W_9_x693 =  23'd823;
localparam signed [DEBIT:0]  W_9_x694 =  23'd833;
localparam signed [DEBIT:0]  W_9_x695 =  23'd907;
localparam signed [DEBIT:0]  W_9_x696 =  23'd954;
localparam signed [DEBIT:0]  W_9_x697 =  23'd952;
localparam signed [DEBIT:0]  W_9_x698 =  23'd950;
localparam signed [DEBIT:0]  W_9_x699 =  23'd959;
localparam signed [DEBIT:0]  W_9_x700 =  23'd970;
localparam signed [DEBIT:0]  W_9_x701 =  23'd967;
localparam signed [DEBIT:0]  W_9_x702 =  23'd960;
localparam signed [DEBIT:0]  W_9_x703 =  23'd961;
localparam signed [DEBIT:0]  W_9_x704 =  23'd953;
localparam signed [DEBIT:0]  W_9_x705 =  23'd918;
localparam signed [DEBIT:0]  W_9_x706 =  23'd881;
localparam signed [DEBIT:0]  W_9_x707 =  23'd792;
localparam signed [DEBIT:0]  W_9_x708 =  23'd722;
localparam signed [DEBIT:0]  W_9_x709 =  23'd621;
localparam signed [DEBIT:0]  W_9_x710 =  23'd522;
localparam signed [DEBIT:0]  W_9_x711 =  23'd473;
localparam signed [DEBIT:0]  W_9_x712 =  23'd458;
localparam signed [DEBIT:0]  W_9_x713 =  23'd469;
localparam signed [DEBIT:0]  W_9_x714 =  23'd437;
localparam signed [DEBIT:0]  W_9_x715 =  23'd450;
localparam signed [DEBIT:0]  W_9_x716 =  23'd485;
localparam signed [DEBIT:0]  W_9_x717 =  23'd607;
localparam signed [DEBIT:0]  W_9_x718 =  23'd752;
localparam signed [DEBIT:0]  W_9_x719 =  23'd821;
localparam signed [DEBIT:0]  W_9_x720 =  23'd929;
localparam signed [DEBIT:0]  W_9_x721 =  23'd1076;
localparam signed [DEBIT:0]  W_9_x722 =  23'd1050;
localparam signed [DEBIT:0]  W_9_x723 =  23'd965;
localparam signed [DEBIT:0]  W_9_x724 =  23'd972;
localparam signed [DEBIT:0]  W_9_x725 =  23'd965;
localparam signed [DEBIT:0]  W_9_x726 =  23'd955;
localparam signed [DEBIT:0]  W_9_x727 =  23'd963;
localparam signed [DEBIT:0]  W_9_x728 =  23'd959;
localparam signed [DEBIT:0]  W_9_x729 =  23'd962;
localparam signed [DEBIT:0]  W_9_x730 =  23'd969;
localparam signed [DEBIT:0]  W_9_x731 =  23'd959;
localparam signed [DEBIT:0]  W_9_x732 =  23'd961;
localparam signed [DEBIT:0]  W_9_x733 =  23'd961;
localparam signed [DEBIT:0]  W_9_x734 =  23'd935;
localparam signed [DEBIT:0]  W_9_x735 =  23'd898;
localparam signed [DEBIT:0]  W_9_x736 =  23'd869;
localparam signed [DEBIT:0]  W_9_x737 =  23'd773;
localparam signed [DEBIT:0]  W_9_x738 =  23'd695;
localparam signed [DEBIT:0]  W_9_x739 =  23'd559;
localparam signed [DEBIT:0]  W_9_x740 =  23'd487;
localparam signed [DEBIT:0]  W_9_x741 =  23'd512;
localparam signed [DEBIT:0]  W_9_x742 =  23'd516;
localparam signed [DEBIT:0]  W_9_x743 =  23'd529;
localparam signed [DEBIT:0]  W_9_x744 =  23'd469;
localparam signed [DEBIT:0]  W_9_x745 =  23'd537;
localparam signed [DEBIT:0]  W_9_x746 =  23'd597;
localparam signed [DEBIT:0]  W_9_x747 =  23'd718;
localparam signed [DEBIT:0]  W_9_x748 =  23'd770;
localparam signed [DEBIT:0]  W_9_x749 =  23'd901;
localparam signed [DEBIT:0]  W_9_x750 =  23'd930;
localparam signed [DEBIT:0]  W_9_x751 =  23'd944;
localparam signed [DEBIT:0]  W_9_x752 =  23'd967;
localparam signed [DEBIT:0]  W_9_x753 =  23'd965;
localparam signed [DEBIT:0]  W_9_x754 =  23'd968;
localparam signed [DEBIT:0]  W_9_x755 =  23'd959;
localparam signed [DEBIT:0]  W_9_x756 =  23'd963;
localparam signed [DEBIT:0]  W_9_x757 =  23'd960;
localparam signed [DEBIT:0]  W_9_x758 =  23'd969;
localparam signed [DEBIT:0]  W_9_x759 =  23'd963;
localparam signed [DEBIT:0]  W_9_x760 =  23'd959;
localparam signed [DEBIT:0]  W_9_x761 =  23'd959;
localparam signed [DEBIT:0]  W_9_x762 =  23'd953;
localparam signed [DEBIT:0]  W_9_x763 =  23'd947;
localparam signed [DEBIT:0]  W_9_x764 =  23'd936;
localparam signed [DEBIT:0]  W_9_x765 =  23'd935;
localparam signed [DEBIT:0]  W_9_x766 =  23'd946;
localparam signed [DEBIT:0]  W_9_x767 =  23'd926;
localparam signed [DEBIT:0]  W_9_x768 =  23'd886;
localparam signed [DEBIT:0]  W_9_x769 =  23'd837;
localparam signed [DEBIT:0]  W_9_x770 =  23'd832;
localparam signed [DEBIT:0]  W_9_x771 =  23'd821;
localparam signed [DEBIT:0]  W_9_x772 =  23'd820;
localparam signed [DEBIT:0]  W_9_x773 =  23'd809;
localparam signed [DEBIT:0]  W_9_x774 =  23'd822;
localparam signed [DEBIT:0]  W_9_x775 =  23'd817;
localparam signed [DEBIT:0]  W_9_x776 =  23'd879;
localparam signed [DEBIT:0]  W_9_x777 =  23'd938;
localparam signed [DEBIT:0]  W_9_x778 =  23'd945;
localparam signed [DEBIT:0]  W_9_x779 =  23'd962;
localparam signed [DEBIT:0]  W_9_x780 =  23'd956;
localparam signed [DEBIT:0]  W_9_x781 =  23'd963;
localparam signed [DEBIT:0]  W_9_x782 =  23'd965;
localparam signed [DEBIT:0]  W_9_x783 =  23'd962;
localparam signed [DEBIT:0]  W_9_x784 =  23'd964;




//****************************    实例化 28*28 共754个实例    *******************************

myram_28X28 #(
.ID(1),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x1),
.W_1(W_1_x1),
.W_2(W_2_x1),
.W_3(W_3_x1),
.W_4(W_4_x1),
.W_5(W_5_x1),
.W_6(W_6_x1),
.W_7(W_7_x1),
.W_8(W_8_x1),
.W_9(W_9_x1)
) u_28X28_x1 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x1),
 .score_0 (score_0_x1),
 .score_1 (score_1_x1),
 .score_2 (score_2_x1),
 .score_3 (score_3_x1),
 .score_4 (score_4_x1),
 .score_5 (score_5_x1),
 .score_6 (score_6_x1),
 .score_7 (score_7_x1),
 .score_8 (score_8_x1),
 .score_9 (score_9_x1)
);
 
myram_28X28 #(
.ID(2),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x2),
.W_1(W_1_x2),
.W_2(W_2_x2),
.W_3(W_3_x2),
.W_4(W_4_x2),
.W_5(W_5_x2),
.W_6(W_6_x2),
.W_7(W_7_x2),
.W_8(W_8_x2),
.W_9(W_9_x2)
) u_28X28_x2 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x2),
 .score_0 (score_0_x2),
 .score_1 (score_1_x2),
 .score_2 (score_2_x2),
 .score_3 (score_3_x2),
 .score_4 (score_4_x2),
 .score_5 (score_5_x2),
 .score_6 (score_6_x2),
 .score_7 (score_7_x2),
 .score_8 (score_8_x2),
 .score_9 (score_9_x2)
);
 
myram_28X28 #(
.ID(3),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x3),
.W_1(W_1_x3),
.W_2(W_2_x3),
.W_3(W_3_x3),
.W_4(W_4_x3),
.W_5(W_5_x3),
.W_6(W_6_x3),
.W_7(W_7_x3),
.W_8(W_8_x3),
.W_9(W_9_x3)
) u_28X28_x3 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x3),
 .score_0 (score_0_x3),
 .score_1 (score_1_x3),
 .score_2 (score_2_x3),
 .score_3 (score_3_x3),
 .score_4 (score_4_x3),
 .score_5 (score_5_x3),
 .score_6 (score_6_x3),
 .score_7 (score_7_x3),
 .score_8 (score_8_x3),
 .score_9 (score_9_x3)
);
 
myram_28X28 #(
.ID(4),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x4),
.W_1(W_1_x4),
.W_2(W_2_x4),
.W_3(W_3_x4),
.W_4(W_4_x4),
.W_5(W_5_x4),
.W_6(W_6_x4),
.W_7(W_7_x4),
.W_8(W_8_x4),
.W_9(W_9_x4)
) u_28X28_x4 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x4),
 .score_0 (score_0_x4),
 .score_1 (score_1_x4),
 .score_2 (score_2_x4),
 .score_3 (score_3_x4),
 .score_4 (score_4_x4),
 .score_5 (score_5_x4),
 .score_6 (score_6_x4),
 .score_7 (score_7_x4),
 .score_8 (score_8_x4),
 .score_9 (score_9_x4)
);
 
myram_28X28 #(
.ID(5),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x5),
.W_1(W_1_x5),
.W_2(W_2_x5),
.W_3(W_3_x5),
.W_4(W_4_x5),
.W_5(W_5_x5),
.W_6(W_6_x5),
.W_7(W_7_x5),
.W_8(W_8_x5),
.W_9(W_9_x5)
) u_28X28_x5 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x5),
 .score_0 (score_0_x5),
 .score_1 (score_1_x5),
 .score_2 (score_2_x5),
 .score_3 (score_3_x5),
 .score_4 (score_4_x5),
 .score_5 (score_5_x5),
 .score_6 (score_6_x5),
 .score_7 (score_7_x5),
 .score_8 (score_8_x5),
 .score_9 (score_9_x5)
);
 
myram_28X28 #(
.ID(6),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x6),
.W_1(W_1_x6),
.W_2(W_2_x6),
.W_3(W_3_x6),
.W_4(W_4_x6),
.W_5(W_5_x6),
.W_6(W_6_x6),
.W_7(W_7_x6),
.W_8(W_8_x6),
.W_9(W_9_x6)
) u_28X28_x6 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x6),
 .score_0 (score_0_x6),
 .score_1 (score_1_x6),
 .score_2 (score_2_x6),
 .score_3 (score_3_x6),
 .score_4 (score_4_x6),
 .score_5 (score_5_x6),
 .score_6 (score_6_x6),
 .score_7 (score_7_x6),
 .score_8 (score_8_x6),
 .score_9 (score_9_x6)
);
 
myram_28X28 #(
.ID(7),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x7),
.W_1(W_1_x7),
.W_2(W_2_x7),
.W_3(W_3_x7),
.W_4(W_4_x7),
.W_5(W_5_x7),
.W_6(W_6_x7),
.W_7(W_7_x7),
.W_8(W_8_x7),
.W_9(W_9_x7)
) u_28X28_x7 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x7),
 .score_0 (score_0_x7),
 .score_1 (score_1_x7),
 .score_2 (score_2_x7),
 .score_3 (score_3_x7),
 .score_4 (score_4_x7),
 .score_5 (score_5_x7),
 .score_6 (score_6_x7),
 .score_7 (score_7_x7),
 .score_8 (score_8_x7),
 .score_9 (score_9_x7)
);
 
myram_28X28 #(
.ID(8),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x8),
.W_1(W_1_x8),
.W_2(W_2_x8),
.W_3(W_3_x8),
.W_4(W_4_x8),
.W_5(W_5_x8),
.W_6(W_6_x8),
.W_7(W_7_x8),
.W_8(W_8_x8),
.W_9(W_9_x8)
) u_28X28_x8 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x8),
 .score_0 (score_0_x8),
 .score_1 (score_1_x8),
 .score_2 (score_2_x8),
 .score_3 (score_3_x8),
 .score_4 (score_4_x8),
 .score_5 (score_5_x8),
 .score_6 (score_6_x8),
 .score_7 (score_7_x8),
 .score_8 (score_8_x8),
 .score_9 (score_9_x8)
);
 
myram_28X28 #(
.ID(9),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x9),
.W_1(W_1_x9),
.W_2(W_2_x9),
.W_3(W_3_x9),
.W_4(W_4_x9),
.W_5(W_5_x9),
.W_6(W_6_x9),
.W_7(W_7_x9),
.W_8(W_8_x9),
.W_9(W_9_x9)
) u_28X28_x9 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x9),
 .score_0 (score_0_x9),
 .score_1 (score_1_x9),
 .score_2 (score_2_x9),
 .score_3 (score_3_x9),
 .score_4 (score_4_x9),
 .score_5 (score_5_x9),
 .score_6 (score_6_x9),
 .score_7 (score_7_x9),
 .score_8 (score_8_x9),
 .score_9 (score_9_x9)
);
 
myram_28X28 #(
.ID(10),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x10),
.W_1(W_1_x10),
.W_2(W_2_x10),
.W_3(W_3_x10),
.W_4(W_4_x10),
.W_5(W_5_x10),
.W_6(W_6_x10),
.W_7(W_7_x10),
.W_8(W_8_x10),
.W_9(W_9_x10)
) u_28X28_x10 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x10),
 .score_0 (score_0_x10),
 .score_1 (score_1_x10),
 .score_2 (score_2_x10),
 .score_3 (score_3_x10),
 .score_4 (score_4_x10),
 .score_5 (score_5_x10),
 .score_6 (score_6_x10),
 .score_7 (score_7_x10),
 .score_8 (score_8_x10),
 .score_9 (score_9_x10)
);
 
myram_28X28 #(
.ID(11),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x11),
.W_1(W_1_x11),
.W_2(W_2_x11),
.W_3(W_3_x11),
.W_4(W_4_x11),
.W_5(W_5_x11),
.W_6(W_6_x11),
.W_7(W_7_x11),
.W_8(W_8_x11),
.W_9(W_9_x11)
) u_28X28_x11 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x11),
 .score_0 (score_0_x11),
 .score_1 (score_1_x11),
 .score_2 (score_2_x11),
 .score_3 (score_3_x11),
 .score_4 (score_4_x11),
 .score_5 (score_5_x11),
 .score_6 (score_6_x11),
 .score_7 (score_7_x11),
 .score_8 (score_8_x11),
 .score_9 (score_9_x11)
);
 
myram_28X28 #(
.ID(12),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x12),
.W_1(W_1_x12),
.W_2(W_2_x12),
.W_3(W_3_x12),
.W_4(W_4_x12),
.W_5(W_5_x12),
.W_6(W_6_x12),
.W_7(W_7_x12),
.W_8(W_8_x12),
.W_9(W_9_x12)
) u_28X28_x12 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x12),
 .score_0 (score_0_x12),
 .score_1 (score_1_x12),
 .score_2 (score_2_x12),
 .score_3 (score_3_x12),
 .score_4 (score_4_x12),
 .score_5 (score_5_x12),
 .score_6 (score_6_x12),
 .score_7 (score_7_x12),
 .score_8 (score_8_x12),
 .score_9 (score_9_x12)
);
 
myram_28X28 #(
.ID(13),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x13),
.W_1(W_1_x13),
.W_2(W_2_x13),
.W_3(W_3_x13),
.W_4(W_4_x13),
.W_5(W_5_x13),
.W_6(W_6_x13),
.W_7(W_7_x13),
.W_8(W_8_x13),
.W_9(W_9_x13)
) u_28X28_x13 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x13),
 .score_0 (score_0_x13),
 .score_1 (score_1_x13),
 .score_2 (score_2_x13),
 .score_3 (score_3_x13),
 .score_4 (score_4_x13),
 .score_5 (score_5_x13),
 .score_6 (score_6_x13),
 .score_7 (score_7_x13),
 .score_8 (score_8_x13),
 .score_9 (score_9_x13)
);
 
myram_28X28 #(
.ID(14),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x14),
.W_1(W_1_x14),
.W_2(W_2_x14),
.W_3(W_3_x14),
.W_4(W_4_x14),
.W_5(W_5_x14),
.W_6(W_6_x14),
.W_7(W_7_x14),
.W_8(W_8_x14),
.W_9(W_9_x14)
) u_28X28_x14 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x14),
 .score_0 (score_0_x14),
 .score_1 (score_1_x14),
 .score_2 (score_2_x14),
 .score_3 (score_3_x14),
 .score_4 (score_4_x14),
 .score_5 (score_5_x14),
 .score_6 (score_6_x14),
 .score_7 (score_7_x14),
 .score_8 (score_8_x14),
 .score_9 (score_9_x14)
);
 
myram_28X28 #(
.ID(15),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x15),
.W_1(W_1_x15),
.W_2(W_2_x15),
.W_3(W_3_x15),
.W_4(W_4_x15),
.W_5(W_5_x15),
.W_6(W_6_x15),
.W_7(W_7_x15),
.W_8(W_8_x15),
.W_9(W_9_x15)
) u_28X28_x15 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x15),
 .score_0 (score_0_x15),
 .score_1 (score_1_x15),
 .score_2 (score_2_x15),
 .score_3 (score_3_x15),
 .score_4 (score_4_x15),
 .score_5 (score_5_x15),
 .score_6 (score_6_x15),
 .score_7 (score_7_x15),
 .score_8 (score_8_x15),
 .score_9 (score_9_x15)
);
 
myram_28X28 #(
.ID(16),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x16),
.W_1(W_1_x16),
.W_2(W_2_x16),
.W_3(W_3_x16),
.W_4(W_4_x16),
.W_5(W_5_x16),
.W_6(W_6_x16),
.W_7(W_7_x16),
.W_8(W_8_x16),
.W_9(W_9_x16)
) u_28X28_x16 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x16),
 .score_0 (score_0_x16),
 .score_1 (score_1_x16),
 .score_2 (score_2_x16),
 .score_3 (score_3_x16),
 .score_4 (score_4_x16),
 .score_5 (score_5_x16),
 .score_6 (score_6_x16),
 .score_7 (score_7_x16),
 .score_8 (score_8_x16),
 .score_9 (score_9_x16)
);
 
myram_28X28 #(
.ID(17),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x17),
.W_1(W_1_x17),
.W_2(W_2_x17),
.W_3(W_3_x17),
.W_4(W_4_x17),
.W_5(W_5_x17),
.W_6(W_6_x17),
.W_7(W_7_x17),
.W_8(W_8_x17),
.W_9(W_9_x17)
) u_28X28_x17 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x17),
 .score_0 (score_0_x17),
 .score_1 (score_1_x17),
 .score_2 (score_2_x17),
 .score_3 (score_3_x17),
 .score_4 (score_4_x17),
 .score_5 (score_5_x17),
 .score_6 (score_6_x17),
 .score_7 (score_7_x17),
 .score_8 (score_8_x17),
 .score_9 (score_9_x17)
);
 
myram_28X28 #(
.ID(18),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x18),
.W_1(W_1_x18),
.W_2(W_2_x18),
.W_3(W_3_x18),
.W_4(W_4_x18),
.W_5(W_5_x18),
.W_6(W_6_x18),
.W_7(W_7_x18),
.W_8(W_8_x18),
.W_9(W_9_x18)
) u_28X28_x18 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x18),
 .score_0 (score_0_x18),
 .score_1 (score_1_x18),
 .score_2 (score_2_x18),
 .score_3 (score_3_x18),
 .score_4 (score_4_x18),
 .score_5 (score_5_x18),
 .score_6 (score_6_x18),
 .score_7 (score_7_x18),
 .score_8 (score_8_x18),
 .score_9 (score_9_x18)
);
 
myram_28X28 #(
.ID(19),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x19),
.W_1(W_1_x19),
.W_2(W_2_x19),
.W_3(W_3_x19),
.W_4(W_4_x19),
.W_5(W_5_x19),
.W_6(W_6_x19),
.W_7(W_7_x19),
.W_8(W_8_x19),
.W_9(W_9_x19)
) u_28X28_x19 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x19),
 .score_0 (score_0_x19),
 .score_1 (score_1_x19),
 .score_2 (score_2_x19),
 .score_3 (score_3_x19),
 .score_4 (score_4_x19),
 .score_5 (score_5_x19),
 .score_6 (score_6_x19),
 .score_7 (score_7_x19),
 .score_8 (score_8_x19),
 .score_9 (score_9_x19)
);
 
myram_28X28 #(
.ID(20),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x20),
.W_1(W_1_x20),
.W_2(W_2_x20),
.W_3(W_3_x20),
.W_4(W_4_x20),
.W_5(W_5_x20),
.W_6(W_6_x20),
.W_7(W_7_x20),
.W_8(W_8_x20),
.W_9(W_9_x20)
) u_28X28_x20 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x20),
 .score_0 (score_0_x20),
 .score_1 (score_1_x20),
 .score_2 (score_2_x20),
 .score_3 (score_3_x20),
 .score_4 (score_4_x20),
 .score_5 (score_5_x20),
 .score_6 (score_6_x20),
 .score_7 (score_7_x20),
 .score_8 (score_8_x20),
 .score_9 (score_9_x20)
);
 
myram_28X28 #(
.ID(21),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x21),
.W_1(W_1_x21),
.W_2(W_2_x21),
.W_3(W_3_x21),
.W_4(W_4_x21),
.W_5(W_5_x21),
.W_6(W_6_x21),
.W_7(W_7_x21),
.W_8(W_8_x21),
.W_9(W_9_x21)
) u_28X28_x21 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x21),
 .score_0 (score_0_x21),
 .score_1 (score_1_x21),
 .score_2 (score_2_x21),
 .score_3 (score_3_x21),
 .score_4 (score_4_x21),
 .score_5 (score_5_x21),
 .score_6 (score_6_x21),
 .score_7 (score_7_x21),
 .score_8 (score_8_x21),
 .score_9 (score_9_x21)
);
 
myram_28X28 #(
.ID(22),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x22),
.W_1(W_1_x22),
.W_2(W_2_x22),
.W_3(W_3_x22),
.W_4(W_4_x22),
.W_5(W_5_x22),
.W_6(W_6_x22),
.W_7(W_7_x22),
.W_8(W_8_x22),
.W_9(W_9_x22)
) u_28X28_x22 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x22),
 .score_0 (score_0_x22),
 .score_1 (score_1_x22),
 .score_2 (score_2_x22),
 .score_3 (score_3_x22),
 .score_4 (score_4_x22),
 .score_5 (score_5_x22),
 .score_6 (score_6_x22),
 .score_7 (score_7_x22),
 .score_8 (score_8_x22),
 .score_9 (score_9_x22)
);
 
myram_28X28 #(
.ID(23),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x23),
.W_1(W_1_x23),
.W_2(W_2_x23),
.W_3(W_3_x23),
.W_4(W_4_x23),
.W_5(W_5_x23),
.W_6(W_6_x23),
.W_7(W_7_x23),
.W_8(W_8_x23),
.W_9(W_9_x23)
) u_28X28_x23 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x23),
 .score_0 (score_0_x23),
 .score_1 (score_1_x23),
 .score_2 (score_2_x23),
 .score_3 (score_3_x23),
 .score_4 (score_4_x23),
 .score_5 (score_5_x23),
 .score_6 (score_6_x23),
 .score_7 (score_7_x23),
 .score_8 (score_8_x23),
 .score_9 (score_9_x23)
);
 
myram_28X28 #(
.ID(24),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x24),
.W_1(W_1_x24),
.W_2(W_2_x24),
.W_3(W_3_x24),
.W_4(W_4_x24),
.W_5(W_5_x24),
.W_6(W_6_x24),
.W_7(W_7_x24),
.W_8(W_8_x24),
.W_9(W_9_x24)
) u_28X28_x24 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x24),
 .score_0 (score_0_x24),
 .score_1 (score_1_x24),
 .score_2 (score_2_x24),
 .score_3 (score_3_x24),
 .score_4 (score_4_x24),
 .score_5 (score_5_x24),
 .score_6 (score_6_x24),
 .score_7 (score_7_x24),
 .score_8 (score_8_x24),
 .score_9 (score_9_x24)
);
 
myram_28X28 #(
.ID(25),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x25),
.W_1(W_1_x25),
.W_2(W_2_x25),
.W_3(W_3_x25),
.W_4(W_4_x25),
.W_5(W_5_x25),
.W_6(W_6_x25),
.W_7(W_7_x25),
.W_8(W_8_x25),
.W_9(W_9_x25)
) u_28X28_x25 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x25),
 .score_0 (score_0_x25),
 .score_1 (score_1_x25),
 .score_2 (score_2_x25),
 .score_3 (score_3_x25),
 .score_4 (score_4_x25),
 .score_5 (score_5_x25),
 .score_6 (score_6_x25),
 .score_7 (score_7_x25),
 .score_8 (score_8_x25),
 .score_9 (score_9_x25)
);
 
myram_28X28 #(
.ID(26),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x26),
.W_1(W_1_x26),
.W_2(W_2_x26),
.W_3(W_3_x26),
.W_4(W_4_x26),
.W_5(W_5_x26),
.W_6(W_6_x26),
.W_7(W_7_x26),
.W_8(W_8_x26),
.W_9(W_9_x26)
) u_28X28_x26 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x26),
 .score_0 (score_0_x26),
 .score_1 (score_1_x26),
 .score_2 (score_2_x26),
 .score_3 (score_3_x26),
 .score_4 (score_4_x26),
 .score_5 (score_5_x26),
 .score_6 (score_6_x26),
 .score_7 (score_7_x26),
 .score_8 (score_8_x26),
 .score_9 (score_9_x26)
);
 
myram_28X28 #(
.ID(27),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x27),
.W_1(W_1_x27),
.W_2(W_2_x27),
.W_3(W_3_x27),
.W_4(W_4_x27),
.W_5(W_5_x27),
.W_6(W_6_x27),
.W_7(W_7_x27),
.W_8(W_8_x27),
.W_9(W_9_x27)
) u_28X28_x27 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x27),
 .score_0 (score_0_x27),
 .score_1 (score_1_x27),
 .score_2 (score_2_x27),
 .score_3 (score_3_x27),
 .score_4 (score_4_x27),
 .score_5 (score_5_x27),
 .score_6 (score_6_x27),
 .score_7 (score_7_x27),
 .score_8 (score_8_x27),
 .score_9 (score_9_x27)
);
 
myram_28X28 #(
.ID(28),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x28),
.W_1(W_1_x28),
.W_2(W_2_x28),
.W_3(W_3_x28),
.W_4(W_4_x28),
.W_5(W_5_x28),
.W_6(W_6_x28),
.W_7(W_7_x28),
.W_8(W_8_x28),
.W_9(W_9_x28)
) u_28X28_x28 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x28),
 .score_0 (score_0_x28),
 .score_1 (score_1_x28),
 .score_2 (score_2_x28),
 .score_3 (score_3_x28),
 .score_4 (score_4_x28),
 .score_5 (score_5_x28),
 .score_6 (score_6_x28),
 .score_7 (score_7_x28),
 .score_8 (score_8_x28),
 .score_9 (score_9_x28)
);
 
myram_28X28 #(
.ID(29),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x29),
.W_1(W_1_x29),
.W_2(W_2_x29),
.W_3(W_3_x29),
.W_4(W_4_x29),
.W_5(W_5_x29),
.W_6(W_6_x29),
.W_7(W_7_x29),
.W_8(W_8_x29),
.W_9(W_9_x29)
) u_28X28_x29 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x29),
 .score_0 (score_0_x29),
 .score_1 (score_1_x29),
 .score_2 (score_2_x29),
 .score_3 (score_3_x29),
 .score_4 (score_4_x29),
 .score_5 (score_5_x29),
 .score_6 (score_6_x29),
 .score_7 (score_7_x29),
 .score_8 (score_8_x29),
 .score_9 (score_9_x29)
);
 
myram_28X28 #(
.ID(30),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x30),
.W_1(W_1_x30),
.W_2(W_2_x30),
.W_3(W_3_x30),
.W_4(W_4_x30),
.W_5(W_5_x30),
.W_6(W_6_x30),
.W_7(W_7_x30),
.W_8(W_8_x30),
.W_9(W_9_x30)
) u_28X28_x30 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x30),
 .score_0 (score_0_x30),
 .score_1 (score_1_x30),
 .score_2 (score_2_x30),
 .score_3 (score_3_x30),
 .score_4 (score_4_x30),
 .score_5 (score_5_x30),
 .score_6 (score_6_x30),
 .score_7 (score_7_x30),
 .score_8 (score_8_x30),
 .score_9 (score_9_x30)
);
 
myram_28X28 #(
.ID(31),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x31),
.W_1(W_1_x31),
.W_2(W_2_x31),
.W_3(W_3_x31),
.W_4(W_4_x31),
.W_5(W_5_x31),
.W_6(W_6_x31),
.W_7(W_7_x31),
.W_8(W_8_x31),
.W_9(W_9_x31)
) u_28X28_x31 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x31),
 .score_0 (score_0_x31),
 .score_1 (score_1_x31),
 .score_2 (score_2_x31),
 .score_3 (score_3_x31),
 .score_4 (score_4_x31),
 .score_5 (score_5_x31),
 .score_6 (score_6_x31),
 .score_7 (score_7_x31),
 .score_8 (score_8_x31),
 .score_9 (score_9_x31)
);
 
myram_28X28 #(
.ID(32),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x32),
.W_1(W_1_x32),
.W_2(W_2_x32),
.W_3(W_3_x32),
.W_4(W_4_x32),
.W_5(W_5_x32),
.W_6(W_6_x32),
.W_7(W_7_x32),
.W_8(W_8_x32),
.W_9(W_9_x32)
) u_28X28_x32 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x32),
 .score_0 (score_0_x32),
 .score_1 (score_1_x32),
 .score_2 (score_2_x32),
 .score_3 (score_3_x32),
 .score_4 (score_4_x32),
 .score_5 (score_5_x32),
 .score_6 (score_6_x32),
 .score_7 (score_7_x32),
 .score_8 (score_8_x32),
 .score_9 (score_9_x32)
);
 
myram_28X28 #(
.ID(33),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x33),
.W_1(W_1_x33),
.W_2(W_2_x33),
.W_3(W_3_x33),
.W_4(W_4_x33),
.W_5(W_5_x33),
.W_6(W_6_x33),
.W_7(W_7_x33),
.W_8(W_8_x33),
.W_9(W_9_x33)
) u_28X28_x33 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x33),
 .score_0 (score_0_x33),
 .score_1 (score_1_x33),
 .score_2 (score_2_x33),
 .score_3 (score_3_x33),
 .score_4 (score_4_x33),
 .score_5 (score_5_x33),
 .score_6 (score_6_x33),
 .score_7 (score_7_x33),
 .score_8 (score_8_x33),
 .score_9 (score_9_x33)
);
 
myram_28X28 #(
.ID(34),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x34),
.W_1(W_1_x34),
.W_2(W_2_x34),
.W_3(W_3_x34),
.W_4(W_4_x34),
.W_5(W_5_x34),
.W_6(W_6_x34),
.W_7(W_7_x34),
.W_8(W_8_x34),
.W_9(W_9_x34)
) u_28X28_x34 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x34),
 .score_0 (score_0_x34),
 .score_1 (score_1_x34),
 .score_2 (score_2_x34),
 .score_3 (score_3_x34),
 .score_4 (score_4_x34),
 .score_5 (score_5_x34),
 .score_6 (score_6_x34),
 .score_7 (score_7_x34),
 .score_8 (score_8_x34),
 .score_9 (score_9_x34)
);
 
myram_28X28 #(
.ID(35),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x35),
.W_1(W_1_x35),
.W_2(W_2_x35),
.W_3(W_3_x35),
.W_4(W_4_x35),
.W_5(W_5_x35),
.W_6(W_6_x35),
.W_7(W_7_x35),
.W_8(W_8_x35),
.W_9(W_9_x35)
) u_28X28_x35 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x35),
 .score_0 (score_0_x35),
 .score_1 (score_1_x35),
 .score_2 (score_2_x35),
 .score_3 (score_3_x35),
 .score_4 (score_4_x35),
 .score_5 (score_5_x35),
 .score_6 (score_6_x35),
 .score_7 (score_7_x35),
 .score_8 (score_8_x35),
 .score_9 (score_9_x35)
);
 
myram_28X28 #(
.ID(36),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x36),
.W_1(W_1_x36),
.W_2(W_2_x36),
.W_3(W_3_x36),
.W_4(W_4_x36),
.W_5(W_5_x36),
.W_6(W_6_x36),
.W_7(W_7_x36),
.W_8(W_8_x36),
.W_9(W_9_x36)
) u_28X28_x36 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x36),
 .score_0 (score_0_x36),
 .score_1 (score_1_x36),
 .score_2 (score_2_x36),
 .score_3 (score_3_x36),
 .score_4 (score_4_x36),
 .score_5 (score_5_x36),
 .score_6 (score_6_x36),
 .score_7 (score_7_x36),
 .score_8 (score_8_x36),
 .score_9 (score_9_x36)
);
 
myram_28X28 #(
.ID(37),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x37),
.W_1(W_1_x37),
.W_2(W_2_x37),
.W_3(W_3_x37),
.W_4(W_4_x37),
.W_5(W_5_x37),
.W_6(W_6_x37),
.W_7(W_7_x37),
.W_8(W_8_x37),
.W_9(W_9_x37)
) u_28X28_x37 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x37),
 .score_0 (score_0_x37),
 .score_1 (score_1_x37),
 .score_2 (score_2_x37),
 .score_3 (score_3_x37),
 .score_4 (score_4_x37),
 .score_5 (score_5_x37),
 .score_6 (score_6_x37),
 .score_7 (score_7_x37),
 .score_8 (score_8_x37),
 .score_9 (score_9_x37)
);
 
myram_28X28 #(
.ID(38),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x38),
.W_1(W_1_x38),
.W_2(W_2_x38),
.W_3(W_3_x38),
.W_4(W_4_x38),
.W_5(W_5_x38),
.W_6(W_6_x38),
.W_7(W_7_x38),
.W_8(W_8_x38),
.W_9(W_9_x38)
) u_28X28_x38 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x38),
 .score_0 (score_0_x38),
 .score_1 (score_1_x38),
 .score_2 (score_2_x38),
 .score_3 (score_3_x38),
 .score_4 (score_4_x38),
 .score_5 (score_5_x38),
 .score_6 (score_6_x38),
 .score_7 (score_7_x38),
 .score_8 (score_8_x38),
 .score_9 (score_9_x38)
);
 
myram_28X28 #(
.ID(39),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x39),
.W_1(W_1_x39),
.W_2(W_2_x39),
.W_3(W_3_x39),
.W_4(W_4_x39),
.W_5(W_5_x39),
.W_6(W_6_x39),
.W_7(W_7_x39),
.W_8(W_8_x39),
.W_9(W_9_x39)
) u_28X28_x39 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x39),
 .score_0 (score_0_x39),
 .score_1 (score_1_x39),
 .score_2 (score_2_x39),
 .score_3 (score_3_x39),
 .score_4 (score_4_x39),
 .score_5 (score_5_x39),
 .score_6 (score_6_x39),
 .score_7 (score_7_x39),
 .score_8 (score_8_x39),
 .score_9 (score_9_x39)
);
 
myram_28X28 #(
.ID(40),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x40),
.W_1(W_1_x40),
.W_2(W_2_x40),
.W_3(W_3_x40),
.W_4(W_4_x40),
.W_5(W_5_x40),
.W_6(W_6_x40),
.W_7(W_7_x40),
.W_8(W_8_x40),
.W_9(W_9_x40)
) u_28X28_x40 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x40),
 .score_0 (score_0_x40),
 .score_1 (score_1_x40),
 .score_2 (score_2_x40),
 .score_3 (score_3_x40),
 .score_4 (score_4_x40),
 .score_5 (score_5_x40),
 .score_6 (score_6_x40),
 .score_7 (score_7_x40),
 .score_8 (score_8_x40),
 .score_9 (score_9_x40)
);
 
myram_28X28 #(
.ID(41),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x41),
.W_1(W_1_x41),
.W_2(W_2_x41),
.W_3(W_3_x41),
.W_4(W_4_x41),
.W_5(W_5_x41),
.W_6(W_6_x41),
.W_7(W_7_x41),
.W_8(W_8_x41),
.W_9(W_9_x41)
) u_28X28_x41 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x41),
 .score_0 (score_0_x41),
 .score_1 (score_1_x41),
 .score_2 (score_2_x41),
 .score_3 (score_3_x41),
 .score_4 (score_4_x41),
 .score_5 (score_5_x41),
 .score_6 (score_6_x41),
 .score_7 (score_7_x41),
 .score_8 (score_8_x41),
 .score_9 (score_9_x41)
);
 
myram_28X28 #(
.ID(42),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x42),
.W_1(W_1_x42),
.W_2(W_2_x42),
.W_3(W_3_x42),
.W_4(W_4_x42),
.W_5(W_5_x42),
.W_6(W_6_x42),
.W_7(W_7_x42),
.W_8(W_8_x42),
.W_9(W_9_x42)
) u_28X28_x42 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x42),
 .score_0 (score_0_x42),
 .score_1 (score_1_x42),
 .score_2 (score_2_x42),
 .score_3 (score_3_x42),
 .score_4 (score_4_x42),
 .score_5 (score_5_x42),
 .score_6 (score_6_x42),
 .score_7 (score_7_x42),
 .score_8 (score_8_x42),
 .score_9 (score_9_x42)
);
 
myram_28X28 #(
.ID(43),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x43),
.W_1(W_1_x43),
.W_2(W_2_x43),
.W_3(W_3_x43),
.W_4(W_4_x43),
.W_5(W_5_x43),
.W_6(W_6_x43),
.W_7(W_7_x43),
.W_8(W_8_x43),
.W_9(W_9_x43)
) u_28X28_x43 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x43),
 .score_0 (score_0_x43),
 .score_1 (score_1_x43),
 .score_2 (score_2_x43),
 .score_3 (score_3_x43),
 .score_4 (score_4_x43),
 .score_5 (score_5_x43),
 .score_6 (score_6_x43),
 .score_7 (score_7_x43),
 .score_8 (score_8_x43),
 .score_9 (score_9_x43)
);
 
myram_28X28 #(
.ID(44),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x44),
.W_1(W_1_x44),
.W_2(W_2_x44),
.W_3(W_3_x44),
.W_4(W_4_x44),
.W_5(W_5_x44),
.W_6(W_6_x44),
.W_7(W_7_x44),
.W_8(W_8_x44),
.W_9(W_9_x44)
) u_28X28_x44 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x44),
 .score_0 (score_0_x44),
 .score_1 (score_1_x44),
 .score_2 (score_2_x44),
 .score_3 (score_3_x44),
 .score_4 (score_4_x44),
 .score_5 (score_5_x44),
 .score_6 (score_6_x44),
 .score_7 (score_7_x44),
 .score_8 (score_8_x44),
 .score_9 (score_9_x44)
);
 
myram_28X28 #(
.ID(45),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x45),
.W_1(W_1_x45),
.W_2(W_2_x45),
.W_3(W_3_x45),
.W_4(W_4_x45),
.W_5(W_5_x45),
.W_6(W_6_x45),
.W_7(W_7_x45),
.W_8(W_8_x45),
.W_9(W_9_x45)
) u_28X28_x45 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x45),
 .score_0 (score_0_x45),
 .score_1 (score_1_x45),
 .score_2 (score_2_x45),
 .score_3 (score_3_x45),
 .score_4 (score_4_x45),
 .score_5 (score_5_x45),
 .score_6 (score_6_x45),
 .score_7 (score_7_x45),
 .score_8 (score_8_x45),
 .score_9 (score_9_x45)
);
 
myram_28X28 #(
.ID(46),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x46),
.W_1(W_1_x46),
.W_2(W_2_x46),
.W_3(W_3_x46),
.W_4(W_4_x46),
.W_5(W_5_x46),
.W_6(W_6_x46),
.W_7(W_7_x46),
.W_8(W_8_x46),
.W_9(W_9_x46)
) u_28X28_x46 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x46),
 .score_0 (score_0_x46),
 .score_1 (score_1_x46),
 .score_2 (score_2_x46),
 .score_3 (score_3_x46),
 .score_4 (score_4_x46),
 .score_5 (score_5_x46),
 .score_6 (score_6_x46),
 .score_7 (score_7_x46),
 .score_8 (score_8_x46),
 .score_9 (score_9_x46)
);
 
myram_28X28 #(
.ID(47),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x47),
.W_1(W_1_x47),
.W_2(W_2_x47),
.W_3(W_3_x47),
.W_4(W_4_x47),
.W_5(W_5_x47),
.W_6(W_6_x47),
.W_7(W_7_x47),
.W_8(W_8_x47),
.W_9(W_9_x47)
) u_28X28_x47 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x47),
 .score_0 (score_0_x47),
 .score_1 (score_1_x47),
 .score_2 (score_2_x47),
 .score_3 (score_3_x47),
 .score_4 (score_4_x47),
 .score_5 (score_5_x47),
 .score_6 (score_6_x47),
 .score_7 (score_7_x47),
 .score_8 (score_8_x47),
 .score_9 (score_9_x47)
);
 
myram_28X28 #(
.ID(48),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x48),
.W_1(W_1_x48),
.W_2(W_2_x48),
.W_3(W_3_x48),
.W_4(W_4_x48),
.W_5(W_5_x48),
.W_6(W_6_x48),
.W_7(W_7_x48),
.W_8(W_8_x48),
.W_9(W_9_x48)
) u_28X28_x48 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x48),
 .score_0 (score_0_x48),
 .score_1 (score_1_x48),
 .score_2 (score_2_x48),
 .score_3 (score_3_x48),
 .score_4 (score_4_x48),
 .score_5 (score_5_x48),
 .score_6 (score_6_x48),
 .score_7 (score_7_x48),
 .score_8 (score_8_x48),
 .score_9 (score_9_x48)
);
 
myram_28X28 #(
.ID(49),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x49),
.W_1(W_1_x49),
.W_2(W_2_x49),
.W_3(W_3_x49),
.W_4(W_4_x49),
.W_5(W_5_x49),
.W_6(W_6_x49),
.W_7(W_7_x49),
.W_8(W_8_x49),
.W_9(W_9_x49)
) u_28X28_x49 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x49),
 .score_0 (score_0_x49),
 .score_1 (score_1_x49),
 .score_2 (score_2_x49),
 .score_3 (score_3_x49),
 .score_4 (score_4_x49),
 .score_5 (score_5_x49),
 .score_6 (score_6_x49),
 .score_7 (score_7_x49),
 .score_8 (score_8_x49),
 .score_9 (score_9_x49)
);
 
myram_28X28 #(
.ID(50),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x50),
.W_1(W_1_x50),
.W_2(W_2_x50),
.W_3(W_3_x50),
.W_4(W_4_x50),
.W_5(W_5_x50),
.W_6(W_6_x50),
.W_7(W_7_x50),
.W_8(W_8_x50),
.W_9(W_9_x50)
) u_28X28_x50 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x50),
 .score_0 (score_0_x50),
 .score_1 (score_1_x50),
 .score_2 (score_2_x50),
 .score_3 (score_3_x50),
 .score_4 (score_4_x50),
 .score_5 (score_5_x50),
 .score_6 (score_6_x50),
 .score_7 (score_7_x50),
 .score_8 (score_8_x50),
 .score_9 (score_9_x50)
);
 
myram_28X28 #(
.ID(51),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x51),
.W_1(W_1_x51),
.W_2(W_2_x51),
.W_3(W_3_x51),
.W_4(W_4_x51),
.W_5(W_5_x51),
.W_6(W_6_x51),
.W_7(W_7_x51),
.W_8(W_8_x51),
.W_9(W_9_x51)
) u_28X28_x51 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x51),
 .score_0 (score_0_x51),
 .score_1 (score_1_x51),
 .score_2 (score_2_x51),
 .score_3 (score_3_x51),
 .score_4 (score_4_x51),
 .score_5 (score_5_x51),
 .score_6 (score_6_x51),
 .score_7 (score_7_x51),
 .score_8 (score_8_x51),
 .score_9 (score_9_x51)
);
 
myram_28X28 #(
.ID(52),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x52),
.W_1(W_1_x52),
.W_2(W_2_x52),
.W_3(W_3_x52),
.W_4(W_4_x52),
.W_5(W_5_x52),
.W_6(W_6_x52),
.W_7(W_7_x52),
.W_8(W_8_x52),
.W_9(W_9_x52)
) u_28X28_x52 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x52),
 .score_0 (score_0_x52),
 .score_1 (score_1_x52),
 .score_2 (score_2_x52),
 .score_3 (score_3_x52),
 .score_4 (score_4_x52),
 .score_5 (score_5_x52),
 .score_6 (score_6_x52),
 .score_7 (score_7_x52),
 .score_8 (score_8_x52),
 .score_9 (score_9_x52)
);
 
myram_28X28 #(
.ID(53),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x53),
.W_1(W_1_x53),
.W_2(W_2_x53),
.W_3(W_3_x53),
.W_4(W_4_x53),
.W_5(W_5_x53),
.W_6(W_6_x53),
.W_7(W_7_x53),
.W_8(W_8_x53),
.W_9(W_9_x53)
) u_28X28_x53 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x53),
 .score_0 (score_0_x53),
 .score_1 (score_1_x53),
 .score_2 (score_2_x53),
 .score_3 (score_3_x53),
 .score_4 (score_4_x53),
 .score_5 (score_5_x53),
 .score_6 (score_6_x53),
 .score_7 (score_7_x53),
 .score_8 (score_8_x53),
 .score_9 (score_9_x53)
);
 
myram_28X28 #(
.ID(54),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x54),
.W_1(W_1_x54),
.W_2(W_2_x54),
.W_3(W_3_x54),
.W_4(W_4_x54),
.W_5(W_5_x54),
.W_6(W_6_x54),
.W_7(W_7_x54),
.W_8(W_8_x54),
.W_9(W_9_x54)
) u_28X28_x54 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x54),
 .score_0 (score_0_x54),
 .score_1 (score_1_x54),
 .score_2 (score_2_x54),
 .score_3 (score_3_x54),
 .score_4 (score_4_x54),
 .score_5 (score_5_x54),
 .score_6 (score_6_x54),
 .score_7 (score_7_x54),
 .score_8 (score_8_x54),
 .score_9 (score_9_x54)
);
 
myram_28X28 #(
.ID(55),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x55),
.W_1(W_1_x55),
.W_2(W_2_x55),
.W_3(W_3_x55),
.W_4(W_4_x55),
.W_5(W_5_x55),
.W_6(W_6_x55),
.W_7(W_7_x55),
.W_8(W_8_x55),
.W_9(W_9_x55)
) u_28X28_x55 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x55),
 .score_0 (score_0_x55),
 .score_1 (score_1_x55),
 .score_2 (score_2_x55),
 .score_3 (score_3_x55),
 .score_4 (score_4_x55),
 .score_5 (score_5_x55),
 .score_6 (score_6_x55),
 .score_7 (score_7_x55),
 .score_8 (score_8_x55),
 .score_9 (score_9_x55)
);
 
myram_28X28 #(
.ID(56),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x56),
.W_1(W_1_x56),
.W_2(W_2_x56),
.W_3(W_3_x56),
.W_4(W_4_x56),
.W_5(W_5_x56),
.W_6(W_6_x56),
.W_7(W_7_x56),
.W_8(W_8_x56),
.W_9(W_9_x56)
) u_28X28_x56 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x56),
 .score_0 (score_0_x56),
 .score_1 (score_1_x56),
 .score_2 (score_2_x56),
 .score_3 (score_3_x56),
 .score_4 (score_4_x56),
 .score_5 (score_5_x56),
 .score_6 (score_6_x56),
 .score_7 (score_7_x56),
 .score_8 (score_8_x56),
 .score_9 (score_9_x56)
);
 
myram_28X28 #(
.ID(57),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x57),
.W_1(W_1_x57),
.W_2(W_2_x57),
.W_3(W_3_x57),
.W_4(W_4_x57),
.W_5(W_5_x57),
.W_6(W_6_x57),
.W_7(W_7_x57),
.W_8(W_8_x57),
.W_9(W_9_x57)
) u_28X28_x57 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x57),
 .score_0 (score_0_x57),
 .score_1 (score_1_x57),
 .score_2 (score_2_x57),
 .score_3 (score_3_x57),
 .score_4 (score_4_x57),
 .score_5 (score_5_x57),
 .score_6 (score_6_x57),
 .score_7 (score_7_x57),
 .score_8 (score_8_x57),
 .score_9 (score_9_x57)
);
 
myram_28X28 #(
.ID(58),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x58),
.W_1(W_1_x58),
.W_2(W_2_x58),
.W_3(W_3_x58),
.W_4(W_4_x58),
.W_5(W_5_x58),
.W_6(W_6_x58),
.W_7(W_7_x58),
.W_8(W_8_x58),
.W_9(W_9_x58)
) u_28X28_x58 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x58),
 .score_0 (score_0_x58),
 .score_1 (score_1_x58),
 .score_2 (score_2_x58),
 .score_3 (score_3_x58),
 .score_4 (score_4_x58),
 .score_5 (score_5_x58),
 .score_6 (score_6_x58),
 .score_7 (score_7_x58),
 .score_8 (score_8_x58),
 .score_9 (score_9_x58)
);
 
myram_28X28 #(
.ID(59),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x59),
.W_1(W_1_x59),
.W_2(W_2_x59),
.W_3(W_3_x59),
.W_4(W_4_x59),
.W_5(W_5_x59),
.W_6(W_6_x59),
.W_7(W_7_x59),
.W_8(W_8_x59),
.W_9(W_9_x59)
) u_28X28_x59 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x59),
 .score_0 (score_0_x59),
 .score_1 (score_1_x59),
 .score_2 (score_2_x59),
 .score_3 (score_3_x59),
 .score_4 (score_4_x59),
 .score_5 (score_5_x59),
 .score_6 (score_6_x59),
 .score_7 (score_7_x59),
 .score_8 (score_8_x59),
 .score_9 (score_9_x59)
);
 
myram_28X28 #(
.ID(60),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x60),
.W_1(W_1_x60),
.W_2(W_2_x60),
.W_3(W_3_x60),
.W_4(W_4_x60),
.W_5(W_5_x60),
.W_6(W_6_x60),
.W_7(W_7_x60),
.W_8(W_8_x60),
.W_9(W_9_x60)
) u_28X28_x60 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x60),
 .score_0 (score_0_x60),
 .score_1 (score_1_x60),
 .score_2 (score_2_x60),
 .score_3 (score_3_x60),
 .score_4 (score_4_x60),
 .score_5 (score_5_x60),
 .score_6 (score_6_x60),
 .score_7 (score_7_x60),
 .score_8 (score_8_x60),
 .score_9 (score_9_x60)
);
 
myram_28X28 #(
.ID(61),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x61),
.W_1(W_1_x61),
.W_2(W_2_x61),
.W_3(W_3_x61),
.W_4(W_4_x61),
.W_5(W_5_x61),
.W_6(W_6_x61),
.W_7(W_7_x61),
.W_8(W_8_x61),
.W_9(W_9_x61)
) u_28X28_x61 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x61),
 .score_0 (score_0_x61),
 .score_1 (score_1_x61),
 .score_2 (score_2_x61),
 .score_3 (score_3_x61),
 .score_4 (score_4_x61),
 .score_5 (score_5_x61),
 .score_6 (score_6_x61),
 .score_7 (score_7_x61),
 .score_8 (score_8_x61),
 .score_9 (score_9_x61)
);
 
myram_28X28 #(
.ID(62),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x62),
.W_1(W_1_x62),
.W_2(W_2_x62),
.W_3(W_3_x62),
.W_4(W_4_x62),
.W_5(W_5_x62),
.W_6(W_6_x62),
.W_7(W_7_x62),
.W_8(W_8_x62),
.W_9(W_9_x62)
) u_28X28_x62 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x62),
 .score_0 (score_0_x62),
 .score_1 (score_1_x62),
 .score_2 (score_2_x62),
 .score_3 (score_3_x62),
 .score_4 (score_4_x62),
 .score_5 (score_5_x62),
 .score_6 (score_6_x62),
 .score_7 (score_7_x62),
 .score_8 (score_8_x62),
 .score_9 (score_9_x62)
);
 
myram_28X28 #(
.ID(63),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x63),
.W_1(W_1_x63),
.W_2(W_2_x63),
.W_3(W_3_x63),
.W_4(W_4_x63),
.W_5(W_5_x63),
.W_6(W_6_x63),
.W_7(W_7_x63),
.W_8(W_8_x63),
.W_9(W_9_x63)
) u_28X28_x63 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x63),
 .score_0 (score_0_x63),
 .score_1 (score_1_x63),
 .score_2 (score_2_x63),
 .score_3 (score_3_x63),
 .score_4 (score_4_x63),
 .score_5 (score_5_x63),
 .score_6 (score_6_x63),
 .score_7 (score_7_x63),
 .score_8 (score_8_x63),
 .score_9 (score_9_x63)
);
 
myram_28X28 #(
.ID(64),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x64),
.W_1(W_1_x64),
.W_2(W_2_x64),
.W_3(W_3_x64),
.W_4(W_4_x64),
.W_5(W_5_x64),
.W_6(W_6_x64),
.W_7(W_7_x64),
.W_8(W_8_x64),
.W_9(W_9_x64)
) u_28X28_x64 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x64),
 .score_0 (score_0_x64),
 .score_1 (score_1_x64),
 .score_2 (score_2_x64),
 .score_3 (score_3_x64),
 .score_4 (score_4_x64),
 .score_5 (score_5_x64),
 .score_6 (score_6_x64),
 .score_7 (score_7_x64),
 .score_8 (score_8_x64),
 .score_9 (score_9_x64)
);
 
myram_28X28 #(
.ID(65),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x65),
.W_1(W_1_x65),
.W_2(W_2_x65),
.W_3(W_3_x65),
.W_4(W_4_x65),
.W_5(W_5_x65),
.W_6(W_6_x65),
.W_7(W_7_x65),
.W_8(W_8_x65),
.W_9(W_9_x65)
) u_28X28_x65 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x65),
 .score_0 (score_0_x65),
 .score_1 (score_1_x65),
 .score_2 (score_2_x65),
 .score_3 (score_3_x65),
 .score_4 (score_4_x65),
 .score_5 (score_5_x65),
 .score_6 (score_6_x65),
 .score_7 (score_7_x65),
 .score_8 (score_8_x65),
 .score_9 (score_9_x65)
);
 
myram_28X28 #(
.ID(66),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x66),
.W_1(W_1_x66),
.W_2(W_2_x66),
.W_3(W_3_x66),
.W_4(W_4_x66),
.W_5(W_5_x66),
.W_6(W_6_x66),
.W_7(W_7_x66),
.W_8(W_8_x66),
.W_9(W_9_x66)
) u_28X28_x66 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x66),
 .score_0 (score_0_x66),
 .score_1 (score_1_x66),
 .score_2 (score_2_x66),
 .score_3 (score_3_x66),
 .score_4 (score_4_x66),
 .score_5 (score_5_x66),
 .score_6 (score_6_x66),
 .score_7 (score_7_x66),
 .score_8 (score_8_x66),
 .score_9 (score_9_x66)
);
 
myram_28X28 #(
.ID(67),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x67),
.W_1(W_1_x67),
.W_2(W_2_x67),
.W_3(W_3_x67),
.W_4(W_4_x67),
.W_5(W_5_x67),
.W_6(W_6_x67),
.W_7(W_7_x67),
.W_8(W_8_x67),
.W_9(W_9_x67)
) u_28X28_x67 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x67),
 .score_0 (score_0_x67),
 .score_1 (score_1_x67),
 .score_2 (score_2_x67),
 .score_3 (score_3_x67),
 .score_4 (score_4_x67),
 .score_5 (score_5_x67),
 .score_6 (score_6_x67),
 .score_7 (score_7_x67),
 .score_8 (score_8_x67),
 .score_9 (score_9_x67)
);
 
myram_28X28 #(
.ID(68),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x68),
.W_1(W_1_x68),
.W_2(W_2_x68),
.W_3(W_3_x68),
.W_4(W_4_x68),
.W_5(W_5_x68),
.W_6(W_6_x68),
.W_7(W_7_x68),
.W_8(W_8_x68),
.W_9(W_9_x68)
) u_28X28_x68 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x68),
 .score_0 (score_0_x68),
 .score_1 (score_1_x68),
 .score_2 (score_2_x68),
 .score_3 (score_3_x68),
 .score_4 (score_4_x68),
 .score_5 (score_5_x68),
 .score_6 (score_6_x68),
 .score_7 (score_7_x68),
 .score_8 (score_8_x68),
 .score_9 (score_9_x68)
);
 
myram_28X28 #(
.ID(69),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x69),
.W_1(W_1_x69),
.W_2(W_2_x69),
.W_3(W_3_x69),
.W_4(W_4_x69),
.W_5(W_5_x69),
.W_6(W_6_x69),
.W_7(W_7_x69),
.W_8(W_8_x69),
.W_9(W_9_x69)
) u_28X28_x69 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x69),
 .score_0 (score_0_x69),
 .score_1 (score_1_x69),
 .score_2 (score_2_x69),
 .score_3 (score_3_x69),
 .score_4 (score_4_x69),
 .score_5 (score_5_x69),
 .score_6 (score_6_x69),
 .score_7 (score_7_x69),
 .score_8 (score_8_x69),
 .score_9 (score_9_x69)
);
 
myram_28X28 #(
.ID(70),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x70),
.W_1(W_1_x70),
.W_2(W_2_x70),
.W_3(W_3_x70),
.W_4(W_4_x70),
.W_5(W_5_x70),
.W_6(W_6_x70),
.W_7(W_7_x70),
.W_8(W_8_x70),
.W_9(W_9_x70)
) u_28X28_x70 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x70),
 .score_0 (score_0_x70),
 .score_1 (score_1_x70),
 .score_2 (score_2_x70),
 .score_3 (score_3_x70),
 .score_4 (score_4_x70),
 .score_5 (score_5_x70),
 .score_6 (score_6_x70),
 .score_7 (score_7_x70),
 .score_8 (score_8_x70),
 .score_9 (score_9_x70)
);
 
myram_28X28 #(
.ID(71),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x71),
.W_1(W_1_x71),
.W_2(W_2_x71),
.W_3(W_3_x71),
.W_4(W_4_x71),
.W_5(W_5_x71),
.W_6(W_6_x71),
.W_7(W_7_x71),
.W_8(W_8_x71),
.W_9(W_9_x71)
) u_28X28_x71 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x71),
 .score_0 (score_0_x71),
 .score_1 (score_1_x71),
 .score_2 (score_2_x71),
 .score_3 (score_3_x71),
 .score_4 (score_4_x71),
 .score_5 (score_5_x71),
 .score_6 (score_6_x71),
 .score_7 (score_7_x71),
 .score_8 (score_8_x71),
 .score_9 (score_9_x71)
);
 
myram_28X28 #(
.ID(72),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x72),
.W_1(W_1_x72),
.W_2(W_2_x72),
.W_3(W_3_x72),
.W_4(W_4_x72),
.W_5(W_5_x72),
.W_6(W_6_x72),
.W_7(W_7_x72),
.W_8(W_8_x72),
.W_9(W_9_x72)
) u_28X28_x72 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x72),
 .score_0 (score_0_x72),
 .score_1 (score_1_x72),
 .score_2 (score_2_x72),
 .score_3 (score_3_x72),
 .score_4 (score_4_x72),
 .score_5 (score_5_x72),
 .score_6 (score_6_x72),
 .score_7 (score_7_x72),
 .score_8 (score_8_x72),
 .score_9 (score_9_x72)
);
 
myram_28X28 #(
.ID(73),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x73),
.W_1(W_1_x73),
.W_2(W_2_x73),
.W_3(W_3_x73),
.W_4(W_4_x73),
.W_5(W_5_x73),
.W_6(W_6_x73),
.W_7(W_7_x73),
.W_8(W_8_x73),
.W_9(W_9_x73)
) u_28X28_x73 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x73),
 .score_0 (score_0_x73),
 .score_1 (score_1_x73),
 .score_2 (score_2_x73),
 .score_3 (score_3_x73),
 .score_4 (score_4_x73),
 .score_5 (score_5_x73),
 .score_6 (score_6_x73),
 .score_7 (score_7_x73),
 .score_8 (score_8_x73),
 .score_9 (score_9_x73)
);
 
myram_28X28 #(
.ID(74),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x74),
.W_1(W_1_x74),
.W_2(W_2_x74),
.W_3(W_3_x74),
.W_4(W_4_x74),
.W_5(W_5_x74),
.W_6(W_6_x74),
.W_7(W_7_x74),
.W_8(W_8_x74),
.W_9(W_9_x74)
) u_28X28_x74 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x74),
 .score_0 (score_0_x74),
 .score_1 (score_1_x74),
 .score_2 (score_2_x74),
 .score_3 (score_3_x74),
 .score_4 (score_4_x74),
 .score_5 (score_5_x74),
 .score_6 (score_6_x74),
 .score_7 (score_7_x74),
 .score_8 (score_8_x74),
 .score_9 (score_9_x74)
);
 
myram_28X28 #(
.ID(75),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x75),
.W_1(W_1_x75),
.W_2(W_2_x75),
.W_3(W_3_x75),
.W_4(W_4_x75),
.W_5(W_5_x75),
.W_6(W_6_x75),
.W_7(W_7_x75),
.W_8(W_8_x75),
.W_9(W_9_x75)
) u_28X28_x75 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x75),
 .score_0 (score_0_x75),
 .score_1 (score_1_x75),
 .score_2 (score_2_x75),
 .score_3 (score_3_x75),
 .score_4 (score_4_x75),
 .score_5 (score_5_x75),
 .score_6 (score_6_x75),
 .score_7 (score_7_x75),
 .score_8 (score_8_x75),
 .score_9 (score_9_x75)
);
 
myram_28X28 #(
.ID(76),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x76),
.W_1(W_1_x76),
.W_2(W_2_x76),
.W_3(W_3_x76),
.W_4(W_4_x76),
.W_5(W_5_x76),
.W_6(W_6_x76),
.W_7(W_7_x76),
.W_8(W_8_x76),
.W_9(W_9_x76)
) u_28X28_x76 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x76),
 .score_0 (score_0_x76),
 .score_1 (score_1_x76),
 .score_2 (score_2_x76),
 .score_3 (score_3_x76),
 .score_4 (score_4_x76),
 .score_5 (score_5_x76),
 .score_6 (score_6_x76),
 .score_7 (score_7_x76),
 .score_8 (score_8_x76),
 .score_9 (score_9_x76)
);
 
myram_28X28 #(
.ID(77),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x77),
.W_1(W_1_x77),
.W_2(W_2_x77),
.W_3(W_3_x77),
.W_4(W_4_x77),
.W_5(W_5_x77),
.W_6(W_6_x77),
.W_7(W_7_x77),
.W_8(W_8_x77),
.W_9(W_9_x77)
) u_28X28_x77 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x77),
 .score_0 (score_0_x77),
 .score_1 (score_1_x77),
 .score_2 (score_2_x77),
 .score_3 (score_3_x77),
 .score_4 (score_4_x77),
 .score_5 (score_5_x77),
 .score_6 (score_6_x77),
 .score_7 (score_7_x77),
 .score_8 (score_8_x77),
 .score_9 (score_9_x77)
);
 
myram_28X28 #(
.ID(78),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x78),
.W_1(W_1_x78),
.W_2(W_2_x78),
.W_3(W_3_x78),
.W_4(W_4_x78),
.W_5(W_5_x78),
.W_6(W_6_x78),
.W_7(W_7_x78),
.W_8(W_8_x78),
.W_9(W_9_x78)
) u_28X28_x78 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x78),
 .score_0 (score_0_x78),
 .score_1 (score_1_x78),
 .score_2 (score_2_x78),
 .score_3 (score_3_x78),
 .score_4 (score_4_x78),
 .score_5 (score_5_x78),
 .score_6 (score_6_x78),
 .score_7 (score_7_x78),
 .score_8 (score_8_x78),
 .score_9 (score_9_x78)
);
 
myram_28X28 #(
.ID(79),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x79),
.W_1(W_1_x79),
.W_2(W_2_x79),
.W_3(W_3_x79),
.W_4(W_4_x79),
.W_5(W_5_x79),
.W_6(W_6_x79),
.W_7(W_7_x79),
.W_8(W_8_x79),
.W_9(W_9_x79)
) u_28X28_x79 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x79),
 .score_0 (score_0_x79),
 .score_1 (score_1_x79),
 .score_2 (score_2_x79),
 .score_3 (score_3_x79),
 .score_4 (score_4_x79),
 .score_5 (score_5_x79),
 .score_6 (score_6_x79),
 .score_7 (score_7_x79),
 .score_8 (score_8_x79),
 .score_9 (score_9_x79)
);
 
myram_28X28 #(
.ID(80),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x80),
.W_1(W_1_x80),
.W_2(W_2_x80),
.W_3(W_3_x80),
.W_4(W_4_x80),
.W_5(W_5_x80),
.W_6(W_6_x80),
.W_7(W_7_x80),
.W_8(W_8_x80),
.W_9(W_9_x80)
) u_28X28_x80 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x80),
 .score_0 (score_0_x80),
 .score_1 (score_1_x80),
 .score_2 (score_2_x80),
 .score_3 (score_3_x80),
 .score_4 (score_4_x80),
 .score_5 (score_5_x80),
 .score_6 (score_6_x80),
 .score_7 (score_7_x80),
 .score_8 (score_8_x80),
 .score_9 (score_9_x80)
);
 
myram_28X28 #(
.ID(81),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x81),
.W_1(W_1_x81),
.W_2(W_2_x81),
.W_3(W_3_x81),
.W_4(W_4_x81),
.W_5(W_5_x81),
.W_6(W_6_x81),
.W_7(W_7_x81),
.W_8(W_8_x81),
.W_9(W_9_x81)
) u_28X28_x81 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x81),
 .score_0 (score_0_x81),
 .score_1 (score_1_x81),
 .score_2 (score_2_x81),
 .score_3 (score_3_x81),
 .score_4 (score_4_x81),
 .score_5 (score_5_x81),
 .score_6 (score_6_x81),
 .score_7 (score_7_x81),
 .score_8 (score_8_x81),
 .score_9 (score_9_x81)
);
 
myram_28X28 #(
.ID(82),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x82),
.W_1(W_1_x82),
.W_2(W_2_x82),
.W_3(W_3_x82),
.W_4(W_4_x82),
.W_5(W_5_x82),
.W_6(W_6_x82),
.W_7(W_7_x82),
.W_8(W_8_x82),
.W_9(W_9_x82)
) u_28X28_x82 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x82),
 .score_0 (score_0_x82),
 .score_1 (score_1_x82),
 .score_2 (score_2_x82),
 .score_3 (score_3_x82),
 .score_4 (score_4_x82),
 .score_5 (score_5_x82),
 .score_6 (score_6_x82),
 .score_7 (score_7_x82),
 .score_8 (score_8_x82),
 .score_9 (score_9_x82)
);
 
myram_28X28 #(
.ID(83),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x83),
.W_1(W_1_x83),
.W_2(W_2_x83),
.W_3(W_3_x83),
.W_4(W_4_x83),
.W_5(W_5_x83),
.W_6(W_6_x83),
.W_7(W_7_x83),
.W_8(W_8_x83),
.W_9(W_9_x83)
) u_28X28_x83 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x83),
 .score_0 (score_0_x83),
 .score_1 (score_1_x83),
 .score_2 (score_2_x83),
 .score_3 (score_3_x83),
 .score_4 (score_4_x83),
 .score_5 (score_5_x83),
 .score_6 (score_6_x83),
 .score_7 (score_7_x83),
 .score_8 (score_8_x83),
 .score_9 (score_9_x83)
);
 
myram_28X28 #(
.ID(84),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x84),
.W_1(W_1_x84),
.W_2(W_2_x84),
.W_3(W_3_x84),
.W_4(W_4_x84),
.W_5(W_5_x84),
.W_6(W_6_x84),
.W_7(W_7_x84),
.W_8(W_8_x84),
.W_9(W_9_x84)
) u_28X28_x84 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x84),
 .score_0 (score_0_x84),
 .score_1 (score_1_x84),
 .score_2 (score_2_x84),
 .score_3 (score_3_x84),
 .score_4 (score_4_x84),
 .score_5 (score_5_x84),
 .score_6 (score_6_x84),
 .score_7 (score_7_x84),
 .score_8 (score_8_x84),
 .score_9 (score_9_x84)
);
 
myram_28X28 #(
.ID(85),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x85),
.W_1(W_1_x85),
.W_2(W_2_x85),
.W_3(W_3_x85),
.W_4(W_4_x85),
.W_5(W_5_x85),
.W_6(W_6_x85),
.W_7(W_7_x85),
.W_8(W_8_x85),
.W_9(W_9_x85)
) u_28X28_x85 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x85),
 .score_0 (score_0_x85),
 .score_1 (score_1_x85),
 .score_2 (score_2_x85),
 .score_3 (score_3_x85),
 .score_4 (score_4_x85),
 .score_5 (score_5_x85),
 .score_6 (score_6_x85),
 .score_7 (score_7_x85),
 .score_8 (score_8_x85),
 .score_9 (score_9_x85)
);
 
myram_28X28 #(
.ID(86),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x86),
.W_1(W_1_x86),
.W_2(W_2_x86),
.W_3(W_3_x86),
.W_4(W_4_x86),
.W_5(W_5_x86),
.W_6(W_6_x86),
.W_7(W_7_x86),
.W_8(W_8_x86),
.W_9(W_9_x86)
) u_28X28_x86 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x86),
 .score_0 (score_0_x86),
 .score_1 (score_1_x86),
 .score_2 (score_2_x86),
 .score_3 (score_3_x86),
 .score_4 (score_4_x86),
 .score_5 (score_5_x86),
 .score_6 (score_6_x86),
 .score_7 (score_7_x86),
 .score_8 (score_8_x86),
 .score_9 (score_9_x86)
);
 
myram_28X28 #(
.ID(87),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x87),
.W_1(W_1_x87),
.W_2(W_2_x87),
.W_3(W_3_x87),
.W_4(W_4_x87),
.W_5(W_5_x87),
.W_6(W_6_x87),
.W_7(W_7_x87),
.W_8(W_8_x87),
.W_9(W_9_x87)
) u_28X28_x87 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x87),
 .score_0 (score_0_x87),
 .score_1 (score_1_x87),
 .score_2 (score_2_x87),
 .score_3 (score_3_x87),
 .score_4 (score_4_x87),
 .score_5 (score_5_x87),
 .score_6 (score_6_x87),
 .score_7 (score_7_x87),
 .score_8 (score_8_x87),
 .score_9 (score_9_x87)
);
 
myram_28X28 #(
.ID(88),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x88),
.W_1(W_1_x88),
.W_2(W_2_x88),
.W_3(W_3_x88),
.W_4(W_4_x88),
.W_5(W_5_x88),
.W_6(W_6_x88),
.W_7(W_7_x88),
.W_8(W_8_x88),
.W_9(W_9_x88)
) u_28X28_x88 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x88),
 .score_0 (score_0_x88),
 .score_1 (score_1_x88),
 .score_2 (score_2_x88),
 .score_3 (score_3_x88),
 .score_4 (score_4_x88),
 .score_5 (score_5_x88),
 .score_6 (score_6_x88),
 .score_7 (score_7_x88),
 .score_8 (score_8_x88),
 .score_9 (score_9_x88)
);
 
myram_28X28 #(
.ID(89),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x89),
.W_1(W_1_x89),
.W_2(W_2_x89),
.W_3(W_3_x89),
.W_4(W_4_x89),
.W_5(W_5_x89),
.W_6(W_6_x89),
.W_7(W_7_x89),
.W_8(W_8_x89),
.W_9(W_9_x89)
) u_28X28_x89 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x89),
 .score_0 (score_0_x89),
 .score_1 (score_1_x89),
 .score_2 (score_2_x89),
 .score_3 (score_3_x89),
 .score_4 (score_4_x89),
 .score_5 (score_5_x89),
 .score_6 (score_6_x89),
 .score_7 (score_7_x89),
 .score_8 (score_8_x89),
 .score_9 (score_9_x89)
);
 
myram_28X28 #(
.ID(90),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x90),
.W_1(W_1_x90),
.W_2(W_2_x90),
.W_3(W_3_x90),
.W_4(W_4_x90),
.W_5(W_5_x90),
.W_6(W_6_x90),
.W_7(W_7_x90),
.W_8(W_8_x90),
.W_9(W_9_x90)
) u_28X28_x90 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x90),
 .score_0 (score_0_x90),
 .score_1 (score_1_x90),
 .score_2 (score_2_x90),
 .score_3 (score_3_x90),
 .score_4 (score_4_x90),
 .score_5 (score_5_x90),
 .score_6 (score_6_x90),
 .score_7 (score_7_x90),
 .score_8 (score_8_x90),
 .score_9 (score_9_x90)
);
 
myram_28X28 #(
.ID(91),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x91),
.W_1(W_1_x91),
.W_2(W_2_x91),
.W_3(W_3_x91),
.W_4(W_4_x91),
.W_5(W_5_x91),
.W_6(W_6_x91),
.W_7(W_7_x91),
.W_8(W_8_x91),
.W_9(W_9_x91)
) u_28X28_x91 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x91),
 .score_0 (score_0_x91),
 .score_1 (score_1_x91),
 .score_2 (score_2_x91),
 .score_3 (score_3_x91),
 .score_4 (score_4_x91),
 .score_5 (score_5_x91),
 .score_6 (score_6_x91),
 .score_7 (score_7_x91),
 .score_8 (score_8_x91),
 .score_9 (score_9_x91)
);
 
myram_28X28 #(
.ID(92),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x92),
.W_1(W_1_x92),
.W_2(W_2_x92),
.W_3(W_3_x92),
.W_4(W_4_x92),
.W_5(W_5_x92),
.W_6(W_6_x92),
.W_7(W_7_x92),
.W_8(W_8_x92),
.W_9(W_9_x92)
) u_28X28_x92 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x92),
 .score_0 (score_0_x92),
 .score_1 (score_1_x92),
 .score_2 (score_2_x92),
 .score_3 (score_3_x92),
 .score_4 (score_4_x92),
 .score_5 (score_5_x92),
 .score_6 (score_6_x92),
 .score_7 (score_7_x92),
 .score_8 (score_8_x92),
 .score_9 (score_9_x92)
);
 
myram_28X28 #(
.ID(93),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x93),
.W_1(W_1_x93),
.W_2(W_2_x93),
.W_3(W_3_x93),
.W_4(W_4_x93),
.W_5(W_5_x93),
.W_6(W_6_x93),
.W_7(W_7_x93),
.W_8(W_8_x93),
.W_9(W_9_x93)
) u_28X28_x93 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x93),
 .score_0 (score_0_x93),
 .score_1 (score_1_x93),
 .score_2 (score_2_x93),
 .score_3 (score_3_x93),
 .score_4 (score_4_x93),
 .score_5 (score_5_x93),
 .score_6 (score_6_x93),
 .score_7 (score_7_x93),
 .score_8 (score_8_x93),
 .score_9 (score_9_x93)
);
 
myram_28X28 #(
.ID(94),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x94),
.W_1(W_1_x94),
.W_2(W_2_x94),
.W_3(W_3_x94),
.W_4(W_4_x94),
.W_5(W_5_x94),
.W_6(W_6_x94),
.W_7(W_7_x94),
.W_8(W_8_x94),
.W_9(W_9_x94)
) u_28X28_x94 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x94),
 .score_0 (score_0_x94),
 .score_1 (score_1_x94),
 .score_2 (score_2_x94),
 .score_3 (score_3_x94),
 .score_4 (score_4_x94),
 .score_5 (score_5_x94),
 .score_6 (score_6_x94),
 .score_7 (score_7_x94),
 .score_8 (score_8_x94),
 .score_9 (score_9_x94)
);
 
myram_28X28 #(
.ID(95),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x95),
.W_1(W_1_x95),
.W_2(W_2_x95),
.W_3(W_3_x95),
.W_4(W_4_x95),
.W_5(W_5_x95),
.W_6(W_6_x95),
.W_7(W_7_x95),
.W_8(W_8_x95),
.W_9(W_9_x95)
) u_28X28_x95 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x95),
 .score_0 (score_0_x95),
 .score_1 (score_1_x95),
 .score_2 (score_2_x95),
 .score_3 (score_3_x95),
 .score_4 (score_4_x95),
 .score_5 (score_5_x95),
 .score_6 (score_6_x95),
 .score_7 (score_7_x95),
 .score_8 (score_8_x95),
 .score_9 (score_9_x95)
);
 
myram_28X28 #(
.ID(96),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x96),
.W_1(W_1_x96),
.W_2(W_2_x96),
.W_3(W_3_x96),
.W_4(W_4_x96),
.W_5(W_5_x96),
.W_6(W_6_x96),
.W_7(W_7_x96),
.W_8(W_8_x96),
.W_9(W_9_x96)
) u_28X28_x96 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x96),
 .score_0 (score_0_x96),
 .score_1 (score_1_x96),
 .score_2 (score_2_x96),
 .score_3 (score_3_x96),
 .score_4 (score_4_x96),
 .score_5 (score_5_x96),
 .score_6 (score_6_x96),
 .score_7 (score_7_x96),
 .score_8 (score_8_x96),
 .score_9 (score_9_x96)
);
 
myram_28X28 #(
.ID(97),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x97),
.W_1(W_1_x97),
.W_2(W_2_x97),
.W_3(W_3_x97),
.W_4(W_4_x97),
.W_5(W_5_x97),
.W_6(W_6_x97),
.W_7(W_7_x97),
.W_8(W_8_x97),
.W_9(W_9_x97)
) u_28X28_x97 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x97),
 .score_0 (score_0_x97),
 .score_1 (score_1_x97),
 .score_2 (score_2_x97),
 .score_3 (score_3_x97),
 .score_4 (score_4_x97),
 .score_5 (score_5_x97),
 .score_6 (score_6_x97),
 .score_7 (score_7_x97),
 .score_8 (score_8_x97),
 .score_9 (score_9_x97)
);
 
myram_28X28 #(
.ID(98),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x98),
.W_1(W_1_x98),
.W_2(W_2_x98),
.W_3(W_3_x98),
.W_4(W_4_x98),
.W_5(W_5_x98),
.W_6(W_6_x98),
.W_7(W_7_x98),
.W_8(W_8_x98),
.W_9(W_9_x98)
) u_28X28_x98 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x98),
 .score_0 (score_0_x98),
 .score_1 (score_1_x98),
 .score_2 (score_2_x98),
 .score_3 (score_3_x98),
 .score_4 (score_4_x98),
 .score_5 (score_5_x98),
 .score_6 (score_6_x98),
 .score_7 (score_7_x98),
 .score_8 (score_8_x98),
 .score_9 (score_9_x98)
);
 
myram_28X28 #(
.ID(99),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x99),
.W_1(W_1_x99),
.W_2(W_2_x99),
.W_3(W_3_x99),
.W_4(W_4_x99),
.W_5(W_5_x99),
.W_6(W_6_x99),
.W_7(W_7_x99),
.W_8(W_8_x99),
.W_9(W_9_x99)
) u_28X28_x99 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x99),
 .score_0 (score_0_x99),
 .score_1 (score_1_x99),
 .score_2 (score_2_x99),
 .score_3 (score_3_x99),
 .score_4 (score_4_x99),
 .score_5 (score_5_x99),
 .score_6 (score_6_x99),
 .score_7 (score_7_x99),
 .score_8 (score_8_x99),
 .score_9 (score_9_x99)
);
 
myram_28X28 #(
.ID(100),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x100),
.W_1(W_1_x100),
.W_2(W_2_x100),
.W_3(W_3_x100),
.W_4(W_4_x100),
.W_5(W_5_x100),
.W_6(W_6_x100),
.W_7(W_7_x100),
.W_8(W_8_x100),
.W_9(W_9_x100)
) u_28X28_x100 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x100),
 .score_0 (score_0_x100),
 .score_1 (score_1_x100),
 .score_2 (score_2_x100),
 .score_3 (score_3_x100),
 .score_4 (score_4_x100),
 .score_5 (score_5_x100),
 .score_6 (score_6_x100),
 .score_7 (score_7_x100),
 .score_8 (score_8_x100),
 .score_9 (score_9_x100)
);
 
myram_28X28 #(
.ID(101),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x101),
.W_1(W_1_x101),
.W_2(W_2_x101),
.W_3(W_3_x101),
.W_4(W_4_x101),
.W_5(W_5_x101),
.W_6(W_6_x101),
.W_7(W_7_x101),
.W_8(W_8_x101),
.W_9(W_9_x101)
) u_28X28_x101 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x101),
 .score_0 (score_0_x101),
 .score_1 (score_1_x101),
 .score_2 (score_2_x101),
 .score_3 (score_3_x101),
 .score_4 (score_4_x101),
 .score_5 (score_5_x101),
 .score_6 (score_6_x101),
 .score_7 (score_7_x101),
 .score_8 (score_8_x101),
 .score_9 (score_9_x101)
);
 
myram_28X28 #(
.ID(102),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x102),
.W_1(W_1_x102),
.W_2(W_2_x102),
.W_3(W_3_x102),
.W_4(W_4_x102),
.W_5(W_5_x102),
.W_6(W_6_x102),
.W_7(W_7_x102),
.W_8(W_8_x102),
.W_9(W_9_x102)
) u_28X28_x102 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x102),
 .score_0 (score_0_x102),
 .score_1 (score_1_x102),
 .score_2 (score_2_x102),
 .score_3 (score_3_x102),
 .score_4 (score_4_x102),
 .score_5 (score_5_x102),
 .score_6 (score_6_x102),
 .score_7 (score_7_x102),
 .score_8 (score_8_x102),
 .score_9 (score_9_x102)
);
 
myram_28X28 #(
.ID(103),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x103),
.W_1(W_1_x103),
.W_2(W_2_x103),
.W_3(W_3_x103),
.W_4(W_4_x103),
.W_5(W_5_x103),
.W_6(W_6_x103),
.W_7(W_7_x103),
.W_8(W_8_x103),
.W_9(W_9_x103)
) u_28X28_x103 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x103),
 .score_0 (score_0_x103),
 .score_1 (score_1_x103),
 .score_2 (score_2_x103),
 .score_3 (score_3_x103),
 .score_4 (score_4_x103),
 .score_5 (score_5_x103),
 .score_6 (score_6_x103),
 .score_7 (score_7_x103),
 .score_8 (score_8_x103),
 .score_9 (score_9_x103)
);
 
myram_28X28 #(
.ID(104),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x104),
.W_1(W_1_x104),
.W_2(W_2_x104),
.W_3(W_3_x104),
.W_4(W_4_x104),
.W_5(W_5_x104),
.W_6(W_6_x104),
.W_7(W_7_x104),
.W_8(W_8_x104),
.W_9(W_9_x104)
) u_28X28_x104 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x104),
 .score_0 (score_0_x104),
 .score_1 (score_1_x104),
 .score_2 (score_2_x104),
 .score_3 (score_3_x104),
 .score_4 (score_4_x104),
 .score_5 (score_5_x104),
 .score_6 (score_6_x104),
 .score_7 (score_7_x104),
 .score_8 (score_8_x104),
 .score_9 (score_9_x104)
);
 
myram_28X28 #(
.ID(105),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x105),
.W_1(W_1_x105),
.W_2(W_2_x105),
.W_3(W_3_x105),
.W_4(W_4_x105),
.W_5(W_5_x105),
.W_6(W_6_x105),
.W_7(W_7_x105),
.W_8(W_8_x105),
.W_9(W_9_x105)
) u_28X28_x105 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x105),
 .score_0 (score_0_x105),
 .score_1 (score_1_x105),
 .score_2 (score_2_x105),
 .score_3 (score_3_x105),
 .score_4 (score_4_x105),
 .score_5 (score_5_x105),
 .score_6 (score_6_x105),
 .score_7 (score_7_x105),
 .score_8 (score_8_x105),
 .score_9 (score_9_x105)
);
 
myram_28X28 #(
.ID(106),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x106),
.W_1(W_1_x106),
.W_2(W_2_x106),
.W_3(W_3_x106),
.W_4(W_4_x106),
.W_5(W_5_x106),
.W_6(W_6_x106),
.W_7(W_7_x106),
.W_8(W_8_x106),
.W_9(W_9_x106)
) u_28X28_x106 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x106),
 .score_0 (score_0_x106),
 .score_1 (score_1_x106),
 .score_2 (score_2_x106),
 .score_3 (score_3_x106),
 .score_4 (score_4_x106),
 .score_5 (score_5_x106),
 .score_6 (score_6_x106),
 .score_7 (score_7_x106),
 .score_8 (score_8_x106),
 .score_9 (score_9_x106)
);
 
myram_28X28 #(
.ID(107),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x107),
.W_1(W_1_x107),
.W_2(W_2_x107),
.W_3(W_3_x107),
.W_4(W_4_x107),
.W_5(W_5_x107),
.W_6(W_6_x107),
.W_7(W_7_x107),
.W_8(W_8_x107),
.W_9(W_9_x107)
) u_28X28_x107 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x107),
 .score_0 (score_0_x107),
 .score_1 (score_1_x107),
 .score_2 (score_2_x107),
 .score_3 (score_3_x107),
 .score_4 (score_4_x107),
 .score_5 (score_5_x107),
 .score_6 (score_6_x107),
 .score_7 (score_7_x107),
 .score_8 (score_8_x107),
 .score_9 (score_9_x107)
);
 
myram_28X28 #(
.ID(108),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x108),
.W_1(W_1_x108),
.W_2(W_2_x108),
.W_3(W_3_x108),
.W_4(W_4_x108),
.W_5(W_5_x108),
.W_6(W_6_x108),
.W_7(W_7_x108),
.W_8(W_8_x108),
.W_9(W_9_x108)
) u_28X28_x108 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x108),
 .score_0 (score_0_x108),
 .score_1 (score_1_x108),
 .score_2 (score_2_x108),
 .score_3 (score_3_x108),
 .score_4 (score_4_x108),
 .score_5 (score_5_x108),
 .score_6 (score_6_x108),
 .score_7 (score_7_x108),
 .score_8 (score_8_x108),
 .score_9 (score_9_x108)
);
 
myram_28X28 #(
.ID(109),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x109),
.W_1(W_1_x109),
.W_2(W_2_x109),
.W_3(W_3_x109),
.W_4(W_4_x109),
.W_5(W_5_x109),
.W_6(W_6_x109),
.W_7(W_7_x109),
.W_8(W_8_x109),
.W_9(W_9_x109)
) u_28X28_x109 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x109),
 .score_0 (score_0_x109),
 .score_1 (score_1_x109),
 .score_2 (score_2_x109),
 .score_3 (score_3_x109),
 .score_4 (score_4_x109),
 .score_5 (score_5_x109),
 .score_6 (score_6_x109),
 .score_7 (score_7_x109),
 .score_8 (score_8_x109),
 .score_9 (score_9_x109)
);
 
myram_28X28 #(
.ID(110),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x110),
.W_1(W_1_x110),
.W_2(W_2_x110),
.W_3(W_3_x110),
.W_4(W_4_x110),
.W_5(W_5_x110),
.W_6(W_6_x110),
.W_7(W_7_x110),
.W_8(W_8_x110),
.W_9(W_9_x110)
) u_28X28_x110 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x110),
 .score_0 (score_0_x110),
 .score_1 (score_1_x110),
 .score_2 (score_2_x110),
 .score_3 (score_3_x110),
 .score_4 (score_4_x110),
 .score_5 (score_5_x110),
 .score_6 (score_6_x110),
 .score_7 (score_7_x110),
 .score_8 (score_8_x110),
 .score_9 (score_9_x110)
);
 
myram_28X28 #(
.ID(111),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x111),
.W_1(W_1_x111),
.W_2(W_2_x111),
.W_3(W_3_x111),
.W_4(W_4_x111),
.W_5(W_5_x111),
.W_6(W_6_x111),
.W_7(W_7_x111),
.W_8(W_8_x111),
.W_9(W_9_x111)
) u_28X28_x111 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x111),
 .score_0 (score_0_x111),
 .score_1 (score_1_x111),
 .score_2 (score_2_x111),
 .score_3 (score_3_x111),
 .score_4 (score_4_x111),
 .score_5 (score_5_x111),
 .score_6 (score_6_x111),
 .score_7 (score_7_x111),
 .score_8 (score_8_x111),
 .score_9 (score_9_x111)
);
 
myram_28X28 #(
.ID(112),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x112),
.W_1(W_1_x112),
.W_2(W_2_x112),
.W_3(W_3_x112),
.W_4(W_4_x112),
.W_5(W_5_x112),
.W_6(W_6_x112),
.W_7(W_7_x112),
.W_8(W_8_x112),
.W_9(W_9_x112)
) u_28X28_x112 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x112),
 .score_0 (score_0_x112),
 .score_1 (score_1_x112),
 .score_2 (score_2_x112),
 .score_3 (score_3_x112),
 .score_4 (score_4_x112),
 .score_5 (score_5_x112),
 .score_6 (score_6_x112),
 .score_7 (score_7_x112),
 .score_8 (score_8_x112),
 .score_9 (score_9_x112)
);
 
myram_28X28 #(
.ID(113),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x113),
.W_1(W_1_x113),
.W_2(W_2_x113),
.W_3(W_3_x113),
.W_4(W_4_x113),
.W_5(W_5_x113),
.W_6(W_6_x113),
.W_7(W_7_x113),
.W_8(W_8_x113),
.W_9(W_9_x113)
) u_28X28_x113 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x113),
 .score_0 (score_0_x113),
 .score_1 (score_1_x113),
 .score_2 (score_2_x113),
 .score_3 (score_3_x113),
 .score_4 (score_4_x113),
 .score_5 (score_5_x113),
 .score_6 (score_6_x113),
 .score_7 (score_7_x113),
 .score_8 (score_8_x113),
 .score_9 (score_9_x113)
);
 
myram_28X28 #(
.ID(114),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x114),
.W_1(W_1_x114),
.W_2(W_2_x114),
.W_3(W_3_x114),
.W_4(W_4_x114),
.W_5(W_5_x114),
.W_6(W_6_x114),
.W_7(W_7_x114),
.W_8(W_8_x114),
.W_9(W_9_x114)
) u_28X28_x114 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x114),
 .score_0 (score_0_x114),
 .score_1 (score_1_x114),
 .score_2 (score_2_x114),
 .score_3 (score_3_x114),
 .score_4 (score_4_x114),
 .score_5 (score_5_x114),
 .score_6 (score_6_x114),
 .score_7 (score_7_x114),
 .score_8 (score_8_x114),
 .score_9 (score_9_x114)
);
 
myram_28X28 #(
.ID(115),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x115),
.W_1(W_1_x115),
.W_2(W_2_x115),
.W_3(W_3_x115),
.W_4(W_4_x115),
.W_5(W_5_x115),
.W_6(W_6_x115),
.W_7(W_7_x115),
.W_8(W_8_x115),
.W_9(W_9_x115)
) u_28X28_x115 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x115),
 .score_0 (score_0_x115),
 .score_1 (score_1_x115),
 .score_2 (score_2_x115),
 .score_3 (score_3_x115),
 .score_4 (score_4_x115),
 .score_5 (score_5_x115),
 .score_6 (score_6_x115),
 .score_7 (score_7_x115),
 .score_8 (score_8_x115),
 .score_9 (score_9_x115)
);
 
myram_28X28 #(
.ID(116),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x116),
.W_1(W_1_x116),
.W_2(W_2_x116),
.W_3(W_3_x116),
.W_4(W_4_x116),
.W_5(W_5_x116),
.W_6(W_6_x116),
.W_7(W_7_x116),
.W_8(W_8_x116),
.W_9(W_9_x116)
) u_28X28_x116 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x116),
 .score_0 (score_0_x116),
 .score_1 (score_1_x116),
 .score_2 (score_2_x116),
 .score_3 (score_3_x116),
 .score_4 (score_4_x116),
 .score_5 (score_5_x116),
 .score_6 (score_6_x116),
 .score_7 (score_7_x116),
 .score_8 (score_8_x116),
 .score_9 (score_9_x116)
);
 
myram_28X28 #(
.ID(117),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x117),
.W_1(W_1_x117),
.W_2(W_2_x117),
.W_3(W_3_x117),
.W_4(W_4_x117),
.W_5(W_5_x117),
.W_6(W_6_x117),
.W_7(W_7_x117),
.W_8(W_8_x117),
.W_9(W_9_x117)
) u_28X28_x117 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x117),
 .score_0 (score_0_x117),
 .score_1 (score_1_x117),
 .score_2 (score_2_x117),
 .score_3 (score_3_x117),
 .score_4 (score_4_x117),
 .score_5 (score_5_x117),
 .score_6 (score_6_x117),
 .score_7 (score_7_x117),
 .score_8 (score_8_x117),
 .score_9 (score_9_x117)
);
 
myram_28X28 #(
.ID(118),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x118),
.W_1(W_1_x118),
.W_2(W_2_x118),
.W_3(W_3_x118),
.W_4(W_4_x118),
.W_5(W_5_x118),
.W_6(W_6_x118),
.W_7(W_7_x118),
.W_8(W_8_x118),
.W_9(W_9_x118)
) u_28X28_x118 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x118),
 .score_0 (score_0_x118),
 .score_1 (score_1_x118),
 .score_2 (score_2_x118),
 .score_3 (score_3_x118),
 .score_4 (score_4_x118),
 .score_5 (score_5_x118),
 .score_6 (score_6_x118),
 .score_7 (score_7_x118),
 .score_8 (score_8_x118),
 .score_9 (score_9_x118)
);
 
myram_28X28 #(
.ID(119),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x119),
.W_1(W_1_x119),
.W_2(W_2_x119),
.W_3(W_3_x119),
.W_4(W_4_x119),
.W_5(W_5_x119),
.W_6(W_6_x119),
.W_7(W_7_x119),
.W_8(W_8_x119),
.W_9(W_9_x119)
) u_28X28_x119 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x119),
 .score_0 (score_0_x119),
 .score_1 (score_1_x119),
 .score_2 (score_2_x119),
 .score_3 (score_3_x119),
 .score_4 (score_4_x119),
 .score_5 (score_5_x119),
 .score_6 (score_6_x119),
 .score_7 (score_7_x119),
 .score_8 (score_8_x119),
 .score_9 (score_9_x119)
);
 
myram_28X28 #(
.ID(120),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x120),
.W_1(W_1_x120),
.W_2(W_2_x120),
.W_3(W_3_x120),
.W_4(W_4_x120),
.W_5(W_5_x120),
.W_6(W_6_x120),
.W_7(W_7_x120),
.W_8(W_8_x120),
.W_9(W_9_x120)
) u_28X28_x120 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x120),
 .score_0 (score_0_x120),
 .score_1 (score_1_x120),
 .score_2 (score_2_x120),
 .score_3 (score_3_x120),
 .score_4 (score_4_x120),
 .score_5 (score_5_x120),
 .score_6 (score_6_x120),
 .score_7 (score_7_x120),
 .score_8 (score_8_x120),
 .score_9 (score_9_x120)
);
 
myram_28X28 #(
.ID(121),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x121),
.W_1(W_1_x121),
.W_2(W_2_x121),
.W_3(W_3_x121),
.W_4(W_4_x121),
.W_5(W_5_x121),
.W_6(W_6_x121),
.W_7(W_7_x121),
.W_8(W_8_x121),
.W_9(W_9_x121)
) u_28X28_x121 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x121),
 .score_0 (score_0_x121),
 .score_1 (score_1_x121),
 .score_2 (score_2_x121),
 .score_3 (score_3_x121),
 .score_4 (score_4_x121),
 .score_5 (score_5_x121),
 .score_6 (score_6_x121),
 .score_7 (score_7_x121),
 .score_8 (score_8_x121),
 .score_9 (score_9_x121)
);
 
myram_28X28 #(
.ID(122),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x122),
.W_1(W_1_x122),
.W_2(W_2_x122),
.W_3(W_3_x122),
.W_4(W_4_x122),
.W_5(W_5_x122),
.W_6(W_6_x122),
.W_7(W_7_x122),
.W_8(W_8_x122),
.W_9(W_9_x122)
) u_28X28_x122 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x122),
 .score_0 (score_0_x122),
 .score_1 (score_1_x122),
 .score_2 (score_2_x122),
 .score_3 (score_3_x122),
 .score_4 (score_4_x122),
 .score_5 (score_5_x122),
 .score_6 (score_6_x122),
 .score_7 (score_7_x122),
 .score_8 (score_8_x122),
 .score_9 (score_9_x122)
);
 
myram_28X28 #(
.ID(123),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x123),
.W_1(W_1_x123),
.W_2(W_2_x123),
.W_3(W_3_x123),
.W_4(W_4_x123),
.W_5(W_5_x123),
.W_6(W_6_x123),
.W_7(W_7_x123),
.W_8(W_8_x123),
.W_9(W_9_x123)
) u_28X28_x123 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x123),
 .score_0 (score_0_x123),
 .score_1 (score_1_x123),
 .score_2 (score_2_x123),
 .score_3 (score_3_x123),
 .score_4 (score_4_x123),
 .score_5 (score_5_x123),
 .score_6 (score_6_x123),
 .score_7 (score_7_x123),
 .score_8 (score_8_x123),
 .score_9 (score_9_x123)
);
 
myram_28X28 #(
.ID(124),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x124),
.W_1(W_1_x124),
.W_2(W_2_x124),
.W_3(W_3_x124),
.W_4(W_4_x124),
.W_5(W_5_x124),
.W_6(W_6_x124),
.W_7(W_7_x124),
.W_8(W_8_x124),
.W_9(W_9_x124)
) u_28X28_x124 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x124),
 .score_0 (score_0_x124),
 .score_1 (score_1_x124),
 .score_2 (score_2_x124),
 .score_3 (score_3_x124),
 .score_4 (score_4_x124),
 .score_5 (score_5_x124),
 .score_6 (score_6_x124),
 .score_7 (score_7_x124),
 .score_8 (score_8_x124),
 .score_9 (score_9_x124)
);
 
myram_28X28 #(
.ID(125),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x125),
.W_1(W_1_x125),
.W_2(W_2_x125),
.W_3(W_3_x125),
.W_4(W_4_x125),
.W_5(W_5_x125),
.W_6(W_6_x125),
.W_7(W_7_x125),
.W_8(W_8_x125),
.W_9(W_9_x125)
) u_28X28_x125 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x125),
 .score_0 (score_0_x125),
 .score_1 (score_1_x125),
 .score_2 (score_2_x125),
 .score_3 (score_3_x125),
 .score_4 (score_4_x125),
 .score_5 (score_5_x125),
 .score_6 (score_6_x125),
 .score_7 (score_7_x125),
 .score_8 (score_8_x125),
 .score_9 (score_9_x125)
);
 
myram_28X28 #(
.ID(126),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x126),
.W_1(W_1_x126),
.W_2(W_2_x126),
.W_3(W_3_x126),
.W_4(W_4_x126),
.W_5(W_5_x126),
.W_6(W_6_x126),
.W_7(W_7_x126),
.W_8(W_8_x126),
.W_9(W_9_x126)
) u_28X28_x126 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x126),
 .score_0 (score_0_x126),
 .score_1 (score_1_x126),
 .score_2 (score_2_x126),
 .score_3 (score_3_x126),
 .score_4 (score_4_x126),
 .score_5 (score_5_x126),
 .score_6 (score_6_x126),
 .score_7 (score_7_x126),
 .score_8 (score_8_x126),
 .score_9 (score_9_x126)
);
 
myram_28X28 #(
.ID(127),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x127),
.W_1(W_1_x127),
.W_2(W_2_x127),
.W_3(W_3_x127),
.W_4(W_4_x127),
.W_5(W_5_x127),
.W_6(W_6_x127),
.W_7(W_7_x127),
.W_8(W_8_x127),
.W_9(W_9_x127)
) u_28X28_x127 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x127),
 .score_0 (score_0_x127),
 .score_1 (score_1_x127),
 .score_2 (score_2_x127),
 .score_3 (score_3_x127),
 .score_4 (score_4_x127),
 .score_5 (score_5_x127),
 .score_6 (score_6_x127),
 .score_7 (score_7_x127),
 .score_8 (score_8_x127),
 .score_9 (score_9_x127)
);
 
myram_28X28 #(
.ID(128),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x128),
.W_1(W_1_x128),
.W_2(W_2_x128),
.W_3(W_3_x128),
.W_4(W_4_x128),
.W_5(W_5_x128),
.W_6(W_6_x128),
.W_7(W_7_x128),
.W_8(W_8_x128),
.W_9(W_9_x128)
) u_28X28_x128 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x128),
 .score_0 (score_0_x128),
 .score_1 (score_1_x128),
 .score_2 (score_2_x128),
 .score_3 (score_3_x128),
 .score_4 (score_4_x128),
 .score_5 (score_5_x128),
 .score_6 (score_6_x128),
 .score_7 (score_7_x128),
 .score_8 (score_8_x128),
 .score_9 (score_9_x128)
);
 
myram_28X28 #(
.ID(129),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x129),
.W_1(W_1_x129),
.W_2(W_2_x129),
.W_3(W_3_x129),
.W_4(W_4_x129),
.W_5(W_5_x129),
.W_6(W_6_x129),
.W_7(W_7_x129),
.W_8(W_8_x129),
.W_9(W_9_x129)
) u_28X28_x129 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x129),
 .score_0 (score_0_x129),
 .score_1 (score_1_x129),
 .score_2 (score_2_x129),
 .score_3 (score_3_x129),
 .score_4 (score_4_x129),
 .score_5 (score_5_x129),
 .score_6 (score_6_x129),
 .score_7 (score_7_x129),
 .score_8 (score_8_x129),
 .score_9 (score_9_x129)
);
 
myram_28X28 #(
.ID(130),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x130),
.W_1(W_1_x130),
.W_2(W_2_x130),
.W_3(W_3_x130),
.W_4(W_4_x130),
.W_5(W_5_x130),
.W_6(W_6_x130),
.W_7(W_7_x130),
.W_8(W_8_x130),
.W_9(W_9_x130)
) u_28X28_x130 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x130),
 .score_0 (score_0_x130),
 .score_1 (score_1_x130),
 .score_2 (score_2_x130),
 .score_3 (score_3_x130),
 .score_4 (score_4_x130),
 .score_5 (score_5_x130),
 .score_6 (score_6_x130),
 .score_7 (score_7_x130),
 .score_8 (score_8_x130),
 .score_9 (score_9_x130)
);
 
myram_28X28 #(
.ID(131),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x131),
.W_1(W_1_x131),
.W_2(W_2_x131),
.W_3(W_3_x131),
.W_4(W_4_x131),
.W_5(W_5_x131),
.W_6(W_6_x131),
.W_7(W_7_x131),
.W_8(W_8_x131),
.W_9(W_9_x131)
) u_28X28_x131 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x131),
 .score_0 (score_0_x131),
 .score_1 (score_1_x131),
 .score_2 (score_2_x131),
 .score_3 (score_3_x131),
 .score_4 (score_4_x131),
 .score_5 (score_5_x131),
 .score_6 (score_6_x131),
 .score_7 (score_7_x131),
 .score_8 (score_8_x131),
 .score_9 (score_9_x131)
);
 
myram_28X28 #(
.ID(132),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x132),
.W_1(W_1_x132),
.W_2(W_2_x132),
.W_3(W_3_x132),
.W_4(W_4_x132),
.W_5(W_5_x132),
.W_6(W_6_x132),
.W_7(W_7_x132),
.W_8(W_8_x132),
.W_9(W_9_x132)
) u_28X28_x132 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x132),
 .score_0 (score_0_x132),
 .score_1 (score_1_x132),
 .score_2 (score_2_x132),
 .score_3 (score_3_x132),
 .score_4 (score_4_x132),
 .score_5 (score_5_x132),
 .score_6 (score_6_x132),
 .score_7 (score_7_x132),
 .score_8 (score_8_x132),
 .score_9 (score_9_x132)
);
 
myram_28X28 #(
.ID(133),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x133),
.W_1(W_1_x133),
.W_2(W_2_x133),
.W_3(W_3_x133),
.W_4(W_4_x133),
.W_5(W_5_x133),
.W_6(W_6_x133),
.W_7(W_7_x133),
.W_8(W_8_x133),
.W_9(W_9_x133)
) u_28X28_x133 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x133),
 .score_0 (score_0_x133),
 .score_1 (score_1_x133),
 .score_2 (score_2_x133),
 .score_3 (score_3_x133),
 .score_4 (score_4_x133),
 .score_5 (score_5_x133),
 .score_6 (score_6_x133),
 .score_7 (score_7_x133),
 .score_8 (score_8_x133),
 .score_9 (score_9_x133)
);
 
myram_28X28 #(
.ID(134),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x134),
.W_1(W_1_x134),
.W_2(W_2_x134),
.W_3(W_3_x134),
.W_4(W_4_x134),
.W_5(W_5_x134),
.W_6(W_6_x134),
.W_7(W_7_x134),
.W_8(W_8_x134),
.W_9(W_9_x134)
) u_28X28_x134 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x134),
 .score_0 (score_0_x134),
 .score_1 (score_1_x134),
 .score_2 (score_2_x134),
 .score_3 (score_3_x134),
 .score_4 (score_4_x134),
 .score_5 (score_5_x134),
 .score_6 (score_6_x134),
 .score_7 (score_7_x134),
 .score_8 (score_8_x134),
 .score_9 (score_9_x134)
);
 
myram_28X28 #(
.ID(135),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x135),
.W_1(W_1_x135),
.W_2(W_2_x135),
.W_3(W_3_x135),
.W_4(W_4_x135),
.W_5(W_5_x135),
.W_6(W_6_x135),
.W_7(W_7_x135),
.W_8(W_8_x135),
.W_9(W_9_x135)
) u_28X28_x135 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x135),
 .score_0 (score_0_x135),
 .score_1 (score_1_x135),
 .score_2 (score_2_x135),
 .score_3 (score_3_x135),
 .score_4 (score_4_x135),
 .score_5 (score_5_x135),
 .score_6 (score_6_x135),
 .score_7 (score_7_x135),
 .score_8 (score_8_x135),
 .score_9 (score_9_x135)
);
 
myram_28X28 #(
.ID(136),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x136),
.W_1(W_1_x136),
.W_2(W_2_x136),
.W_3(W_3_x136),
.W_4(W_4_x136),
.W_5(W_5_x136),
.W_6(W_6_x136),
.W_7(W_7_x136),
.W_8(W_8_x136),
.W_9(W_9_x136)
) u_28X28_x136 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x136),
 .score_0 (score_0_x136),
 .score_1 (score_1_x136),
 .score_2 (score_2_x136),
 .score_3 (score_3_x136),
 .score_4 (score_4_x136),
 .score_5 (score_5_x136),
 .score_6 (score_6_x136),
 .score_7 (score_7_x136),
 .score_8 (score_8_x136),
 .score_9 (score_9_x136)
);
 
myram_28X28 #(
.ID(137),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x137),
.W_1(W_1_x137),
.W_2(W_2_x137),
.W_3(W_3_x137),
.W_4(W_4_x137),
.W_5(W_5_x137),
.W_6(W_6_x137),
.W_7(W_7_x137),
.W_8(W_8_x137),
.W_9(W_9_x137)
) u_28X28_x137 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x137),
 .score_0 (score_0_x137),
 .score_1 (score_1_x137),
 .score_2 (score_2_x137),
 .score_3 (score_3_x137),
 .score_4 (score_4_x137),
 .score_5 (score_5_x137),
 .score_6 (score_6_x137),
 .score_7 (score_7_x137),
 .score_8 (score_8_x137),
 .score_9 (score_9_x137)
);
 
myram_28X28 #(
.ID(138),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x138),
.W_1(W_1_x138),
.W_2(W_2_x138),
.W_3(W_3_x138),
.W_4(W_4_x138),
.W_5(W_5_x138),
.W_6(W_6_x138),
.W_7(W_7_x138),
.W_8(W_8_x138),
.W_9(W_9_x138)
) u_28X28_x138 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x138),
 .score_0 (score_0_x138),
 .score_1 (score_1_x138),
 .score_2 (score_2_x138),
 .score_3 (score_3_x138),
 .score_4 (score_4_x138),
 .score_5 (score_5_x138),
 .score_6 (score_6_x138),
 .score_7 (score_7_x138),
 .score_8 (score_8_x138),
 .score_9 (score_9_x138)
);
 
myram_28X28 #(
.ID(139),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x139),
.W_1(W_1_x139),
.W_2(W_2_x139),
.W_3(W_3_x139),
.W_4(W_4_x139),
.W_5(W_5_x139),
.W_6(W_6_x139),
.W_7(W_7_x139),
.W_8(W_8_x139),
.W_9(W_9_x139)
) u_28X28_x139 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x139),
 .score_0 (score_0_x139),
 .score_1 (score_1_x139),
 .score_2 (score_2_x139),
 .score_3 (score_3_x139),
 .score_4 (score_4_x139),
 .score_5 (score_5_x139),
 .score_6 (score_6_x139),
 .score_7 (score_7_x139),
 .score_8 (score_8_x139),
 .score_9 (score_9_x139)
);
 
myram_28X28 #(
.ID(140),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x140),
.W_1(W_1_x140),
.W_2(W_2_x140),
.W_3(W_3_x140),
.W_4(W_4_x140),
.W_5(W_5_x140),
.W_6(W_6_x140),
.W_7(W_7_x140),
.W_8(W_8_x140),
.W_9(W_9_x140)
) u_28X28_x140 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x140),
 .score_0 (score_0_x140),
 .score_1 (score_1_x140),
 .score_2 (score_2_x140),
 .score_3 (score_3_x140),
 .score_4 (score_4_x140),
 .score_5 (score_5_x140),
 .score_6 (score_6_x140),
 .score_7 (score_7_x140),
 .score_8 (score_8_x140),
 .score_9 (score_9_x140)
);
 
myram_28X28 #(
.ID(141),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x141),
.W_1(W_1_x141),
.W_2(W_2_x141),
.W_3(W_3_x141),
.W_4(W_4_x141),
.W_5(W_5_x141),
.W_6(W_6_x141),
.W_7(W_7_x141),
.W_8(W_8_x141),
.W_9(W_9_x141)
) u_28X28_x141 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x141),
 .score_0 (score_0_x141),
 .score_1 (score_1_x141),
 .score_2 (score_2_x141),
 .score_3 (score_3_x141),
 .score_4 (score_4_x141),
 .score_5 (score_5_x141),
 .score_6 (score_6_x141),
 .score_7 (score_7_x141),
 .score_8 (score_8_x141),
 .score_9 (score_9_x141)
);
 
myram_28X28 #(
.ID(142),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x142),
.W_1(W_1_x142),
.W_2(W_2_x142),
.W_3(W_3_x142),
.W_4(W_4_x142),
.W_5(W_5_x142),
.W_6(W_6_x142),
.W_7(W_7_x142),
.W_8(W_8_x142),
.W_9(W_9_x142)
) u_28X28_x142 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x142),
 .score_0 (score_0_x142),
 .score_1 (score_1_x142),
 .score_2 (score_2_x142),
 .score_3 (score_3_x142),
 .score_4 (score_4_x142),
 .score_5 (score_5_x142),
 .score_6 (score_6_x142),
 .score_7 (score_7_x142),
 .score_8 (score_8_x142),
 .score_9 (score_9_x142)
);
 
myram_28X28 #(
.ID(143),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x143),
.W_1(W_1_x143),
.W_2(W_2_x143),
.W_3(W_3_x143),
.W_4(W_4_x143),
.W_5(W_5_x143),
.W_6(W_6_x143),
.W_7(W_7_x143),
.W_8(W_8_x143),
.W_9(W_9_x143)
) u_28X28_x143 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x143),
 .score_0 (score_0_x143),
 .score_1 (score_1_x143),
 .score_2 (score_2_x143),
 .score_3 (score_3_x143),
 .score_4 (score_4_x143),
 .score_5 (score_5_x143),
 .score_6 (score_6_x143),
 .score_7 (score_7_x143),
 .score_8 (score_8_x143),
 .score_9 (score_9_x143)
);
 
myram_28X28 #(
.ID(144),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x144),
.W_1(W_1_x144),
.W_2(W_2_x144),
.W_3(W_3_x144),
.W_4(W_4_x144),
.W_5(W_5_x144),
.W_6(W_6_x144),
.W_7(W_7_x144),
.W_8(W_8_x144),
.W_9(W_9_x144)
) u_28X28_x144 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x144),
 .score_0 (score_0_x144),
 .score_1 (score_1_x144),
 .score_2 (score_2_x144),
 .score_3 (score_3_x144),
 .score_4 (score_4_x144),
 .score_5 (score_5_x144),
 .score_6 (score_6_x144),
 .score_7 (score_7_x144),
 .score_8 (score_8_x144),
 .score_9 (score_9_x144)
);
 
myram_28X28 #(
.ID(145),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x145),
.W_1(W_1_x145),
.W_2(W_2_x145),
.W_3(W_3_x145),
.W_4(W_4_x145),
.W_5(W_5_x145),
.W_6(W_6_x145),
.W_7(W_7_x145),
.W_8(W_8_x145),
.W_9(W_9_x145)
) u_28X28_x145 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x145),
 .score_0 (score_0_x145),
 .score_1 (score_1_x145),
 .score_2 (score_2_x145),
 .score_3 (score_3_x145),
 .score_4 (score_4_x145),
 .score_5 (score_5_x145),
 .score_6 (score_6_x145),
 .score_7 (score_7_x145),
 .score_8 (score_8_x145),
 .score_9 (score_9_x145)
);
 
myram_28X28 #(
.ID(146),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x146),
.W_1(W_1_x146),
.W_2(W_2_x146),
.W_3(W_3_x146),
.W_4(W_4_x146),
.W_5(W_5_x146),
.W_6(W_6_x146),
.W_7(W_7_x146),
.W_8(W_8_x146),
.W_9(W_9_x146)
) u_28X28_x146 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x146),
 .score_0 (score_0_x146),
 .score_1 (score_1_x146),
 .score_2 (score_2_x146),
 .score_3 (score_3_x146),
 .score_4 (score_4_x146),
 .score_5 (score_5_x146),
 .score_6 (score_6_x146),
 .score_7 (score_7_x146),
 .score_8 (score_8_x146),
 .score_9 (score_9_x146)
);
 
myram_28X28 #(
.ID(147),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x147),
.W_1(W_1_x147),
.W_2(W_2_x147),
.W_3(W_3_x147),
.W_4(W_4_x147),
.W_5(W_5_x147),
.W_6(W_6_x147),
.W_7(W_7_x147),
.W_8(W_8_x147),
.W_9(W_9_x147)
) u_28X28_x147 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x147),
 .score_0 (score_0_x147),
 .score_1 (score_1_x147),
 .score_2 (score_2_x147),
 .score_3 (score_3_x147),
 .score_4 (score_4_x147),
 .score_5 (score_5_x147),
 .score_6 (score_6_x147),
 .score_7 (score_7_x147),
 .score_8 (score_8_x147),
 .score_9 (score_9_x147)
);
 
myram_28X28 #(
.ID(148),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x148),
.W_1(W_1_x148),
.W_2(W_2_x148),
.W_3(W_3_x148),
.W_4(W_4_x148),
.W_5(W_5_x148),
.W_6(W_6_x148),
.W_7(W_7_x148),
.W_8(W_8_x148),
.W_9(W_9_x148)
) u_28X28_x148 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x148),
 .score_0 (score_0_x148),
 .score_1 (score_1_x148),
 .score_2 (score_2_x148),
 .score_3 (score_3_x148),
 .score_4 (score_4_x148),
 .score_5 (score_5_x148),
 .score_6 (score_6_x148),
 .score_7 (score_7_x148),
 .score_8 (score_8_x148),
 .score_9 (score_9_x148)
);
 
myram_28X28 #(
.ID(149),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x149),
.W_1(W_1_x149),
.W_2(W_2_x149),
.W_3(W_3_x149),
.W_4(W_4_x149),
.W_5(W_5_x149),
.W_6(W_6_x149),
.W_7(W_7_x149),
.W_8(W_8_x149),
.W_9(W_9_x149)
) u_28X28_x149 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x149),
 .score_0 (score_0_x149),
 .score_1 (score_1_x149),
 .score_2 (score_2_x149),
 .score_3 (score_3_x149),
 .score_4 (score_4_x149),
 .score_5 (score_5_x149),
 .score_6 (score_6_x149),
 .score_7 (score_7_x149),
 .score_8 (score_8_x149),
 .score_9 (score_9_x149)
);
 
myram_28X28 #(
.ID(150),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x150),
.W_1(W_1_x150),
.W_2(W_2_x150),
.W_3(W_3_x150),
.W_4(W_4_x150),
.W_5(W_5_x150),
.W_6(W_6_x150),
.W_7(W_7_x150),
.W_8(W_8_x150),
.W_9(W_9_x150)
) u_28X28_x150 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x150),
 .score_0 (score_0_x150),
 .score_1 (score_1_x150),
 .score_2 (score_2_x150),
 .score_3 (score_3_x150),
 .score_4 (score_4_x150),
 .score_5 (score_5_x150),
 .score_6 (score_6_x150),
 .score_7 (score_7_x150),
 .score_8 (score_8_x150),
 .score_9 (score_9_x150)
);
 
myram_28X28 #(
.ID(151),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x151),
.W_1(W_1_x151),
.W_2(W_2_x151),
.W_3(W_3_x151),
.W_4(W_4_x151),
.W_5(W_5_x151),
.W_6(W_6_x151),
.W_7(W_7_x151),
.W_8(W_8_x151),
.W_9(W_9_x151)
) u_28X28_x151 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x151),
 .score_0 (score_0_x151),
 .score_1 (score_1_x151),
 .score_2 (score_2_x151),
 .score_3 (score_3_x151),
 .score_4 (score_4_x151),
 .score_5 (score_5_x151),
 .score_6 (score_6_x151),
 .score_7 (score_7_x151),
 .score_8 (score_8_x151),
 .score_9 (score_9_x151)
);
 
myram_28X28 #(
.ID(152),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x152),
.W_1(W_1_x152),
.W_2(W_2_x152),
.W_3(W_3_x152),
.W_4(W_4_x152),
.W_5(W_5_x152),
.W_6(W_6_x152),
.W_7(W_7_x152),
.W_8(W_8_x152),
.W_9(W_9_x152)
) u_28X28_x152 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x152),
 .score_0 (score_0_x152),
 .score_1 (score_1_x152),
 .score_2 (score_2_x152),
 .score_3 (score_3_x152),
 .score_4 (score_4_x152),
 .score_5 (score_5_x152),
 .score_6 (score_6_x152),
 .score_7 (score_7_x152),
 .score_8 (score_8_x152),
 .score_9 (score_9_x152)
);
 
myram_28X28 #(
.ID(153),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x153),
.W_1(W_1_x153),
.W_2(W_2_x153),
.W_3(W_3_x153),
.W_4(W_4_x153),
.W_5(W_5_x153),
.W_6(W_6_x153),
.W_7(W_7_x153),
.W_8(W_8_x153),
.W_9(W_9_x153)
) u_28X28_x153 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x153),
 .score_0 (score_0_x153),
 .score_1 (score_1_x153),
 .score_2 (score_2_x153),
 .score_3 (score_3_x153),
 .score_4 (score_4_x153),
 .score_5 (score_5_x153),
 .score_6 (score_6_x153),
 .score_7 (score_7_x153),
 .score_8 (score_8_x153),
 .score_9 (score_9_x153)
);
 
myram_28X28 #(
.ID(154),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x154),
.W_1(W_1_x154),
.W_2(W_2_x154),
.W_3(W_3_x154),
.W_4(W_4_x154),
.W_5(W_5_x154),
.W_6(W_6_x154),
.W_7(W_7_x154),
.W_8(W_8_x154),
.W_9(W_9_x154)
) u_28X28_x154 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x154),
 .score_0 (score_0_x154),
 .score_1 (score_1_x154),
 .score_2 (score_2_x154),
 .score_3 (score_3_x154),
 .score_4 (score_4_x154),
 .score_5 (score_5_x154),
 .score_6 (score_6_x154),
 .score_7 (score_7_x154),
 .score_8 (score_8_x154),
 .score_9 (score_9_x154)
);
 
myram_28X28 #(
.ID(155),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x155),
.W_1(W_1_x155),
.W_2(W_2_x155),
.W_3(W_3_x155),
.W_4(W_4_x155),
.W_5(W_5_x155),
.W_6(W_6_x155),
.W_7(W_7_x155),
.W_8(W_8_x155),
.W_9(W_9_x155)
) u_28X28_x155 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x155),
 .score_0 (score_0_x155),
 .score_1 (score_1_x155),
 .score_2 (score_2_x155),
 .score_3 (score_3_x155),
 .score_4 (score_4_x155),
 .score_5 (score_5_x155),
 .score_6 (score_6_x155),
 .score_7 (score_7_x155),
 .score_8 (score_8_x155),
 .score_9 (score_9_x155)
);
 
myram_28X28 #(
.ID(156),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x156),
.W_1(W_1_x156),
.W_2(W_2_x156),
.W_3(W_3_x156),
.W_4(W_4_x156),
.W_5(W_5_x156),
.W_6(W_6_x156),
.W_7(W_7_x156),
.W_8(W_8_x156),
.W_9(W_9_x156)
) u_28X28_x156 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x156),
 .score_0 (score_0_x156),
 .score_1 (score_1_x156),
 .score_2 (score_2_x156),
 .score_3 (score_3_x156),
 .score_4 (score_4_x156),
 .score_5 (score_5_x156),
 .score_6 (score_6_x156),
 .score_7 (score_7_x156),
 .score_8 (score_8_x156),
 .score_9 (score_9_x156)
);
 
myram_28X28 #(
.ID(157),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x157),
.W_1(W_1_x157),
.W_2(W_2_x157),
.W_3(W_3_x157),
.W_4(W_4_x157),
.W_5(W_5_x157),
.W_6(W_6_x157),
.W_7(W_7_x157),
.W_8(W_8_x157),
.W_9(W_9_x157)
) u_28X28_x157 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x157),
 .score_0 (score_0_x157),
 .score_1 (score_1_x157),
 .score_2 (score_2_x157),
 .score_3 (score_3_x157),
 .score_4 (score_4_x157),
 .score_5 (score_5_x157),
 .score_6 (score_6_x157),
 .score_7 (score_7_x157),
 .score_8 (score_8_x157),
 .score_9 (score_9_x157)
);
 
myram_28X28 #(
.ID(158),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x158),
.W_1(W_1_x158),
.W_2(W_2_x158),
.W_3(W_3_x158),
.W_4(W_4_x158),
.W_5(W_5_x158),
.W_6(W_6_x158),
.W_7(W_7_x158),
.W_8(W_8_x158),
.W_9(W_9_x158)
) u_28X28_x158 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x158),
 .score_0 (score_0_x158),
 .score_1 (score_1_x158),
 .score_2 (score_2_x158),
 .score_3 (score_3_x158),
 .score_4 (score_4_x158),
 .score_5 (score_5_x158),
 .score_6 (score_6_x158),
 .score_7 (score_7_x158),
 .score_8 (score_8_x158),
 .score_9 (score_9_x158)
);
 
myram_28X28 #(
.ID(159),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x159),
.W_1(W_1_x159),
.W_2(W_2_x159),
.W_3(W_3_x159),
.W_4(W_4_x159),
.W_5(W_5_x159),
.W_6(W_6_x159),
.W_7(W_7_x159),
.W_8(W_8_x159),
.W_9(W_9_x159)
) u_28X28_x159 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x159),
 .score_0 (score_0_x159),
 .score_1 (score_1_x159),
 .score_2 (score_2_x159),
 .score_3 (score_3_x159),
 .score_4 (score_4_x159),
 .score_5 (score_5_x159),
 .score_6 (score_6_x159),
 .score_7 (score_7_x159),
 .score_8 (score_8_x159),
 .score_9 (score_9_x159)
);
 
myram_28X28 #(
.ID(160),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x160),
.W_1(W_1_x160),
.W_2(W_2_x160),
.W_3(W_3_x160),
.W_4(W_4_x160),
.W_5(W_5_x160),
.W_6(W_6_x160),
.W_7(W_7_x160),
.W_8(W_8_x160),
.W_9(W_9_x160)
) u_28X28_x160 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x160),
 .score_0 (score_0_x160),
 .score_1 (score_1_x160),
 .score_2 (score_2_x160),
 .score_3 (score_3_x160),
 .score_4 (score_4_x160),
 .score_5 (score_5_x160),
 .score_6 (score_6_x160),
 .score_7 (score_7_x160),
 .score_8 (score_8_x160),
 .score_9 (score_9_x160)
);
 
myram_28X28 #(
.ID(161),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x161),
.W_1(W_1_x161),
.W_2(W_2_x161),
.W_3(W_3_x161),
.W_4(W_4_x161),
.W_5(W_5_x161),
.W_6(W_6_x161),
.W_7(W_7_x161),
.W_8(W_8_x161),
.W_9(W_9_x161)
) u_28X28_x161 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x161),
 .score_0 (score_0_x161),
 .score_1 (score_1_x161),
 .score_2 (score_2_x161),
 .score_3 (score_3_x161),
 .score_4 (score_4_x161),
 .score_5 (score_5_x161),
 .score_6 (score_6_x161),
 .score_7 (score_7_x161),
 .score_8 (score_8_x161),
 .score_9 (score_9_x161)
);
 
myram_28X28 #(
.ID(162),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x162),
.W_1(W_1_x162),
.W_2(W_2_x162),
.W_3(W_3_x162),
.W_4(W_4_x162),
.W_5(W_5_x162),
.W_6(W_6_x162),
.W_7(W_7_x162),
.W_8(W_8_x162),
.W_9(W_9_x162)
) u_28X28_x162 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x162),
 .score_0 (score_0_x162),
 .score_1 (score_1_x162),
 .score_2 (score_2_x162),
 .score_3 (score_3_x162),
 .score_4 (score_4_x162),
 .score_5 (score_5_x162),
 .score_6 (score_6_x162),
 .score_7 (score_7_x162),
 .score_8 (score_8_x162),
 .score_9 (score_9_x162)
);
 
myram_28X28 #(
.ID(163),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x163),
.W_1(W_1_x163),
.W_2(W_2_x163),
.W_3(W_3_x163),
.W_4(W_4_x163),
.W_5(W_5_x163),
.W_6(W_6_x163),
.W_7(W_7_x163),
.W_8(W_8_x163),
.W_9(W_9_x163)
) u_28X28_x163 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x163),
 .score_0 (score_0_x163),
 .score_1 (score_1_x163),
 .score_2 (score_2_x163),
 .score_3 (score_3_x163),
 .score_4 (score_4_x163),
 .score_5 (score_5_x163),
 .score_6 (score_6_x163),
 .score_7 (score_7_x163),
 .score_8 (score_8_x163),
 .score_9 (score_9_x163)
);
 
myram_28X28 #(
.ID(164),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x164),
.W_1(W_1_x164),
.W_2(W_2_x164),
.W_3(W_3_x164),
.W_4(W_4_x164),
.W_5(W_5_x164),
.W_6(W_6_x164),
.W_7(W_7_x164),
.W_8(W_8_x164),
.W_9(W_9_x164)
) u_28X28_x164 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x164),
 .score_0 (score_0_x164),
 .score_1 (score_1_x164),
 .score_2 (score_2_x164),
 .score_3 (score_3_x164),
 .score_4 (score_4_x164),
 .score_5 (score_5_x164),
 .score_6 (score_6_x164),
 .score_7 (score_7_x164),
 .score_8 (score_8_x164),
 .score_9 (score_9_x164)
);
 
myram_28X28 #(
.ID(165),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x165),
.W_1(W_1_x165),
.W_2(W_2_x165),
.W_3(W_3_x165),
.W_4(W_4_x165),
.W_5(W_5_x165),
.W_6(W_6_x165),
.W_7(W_7_x165),
.W_8(W_8_x165),
.W_9(W_9_x165)
) u_28X28_x165 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x165),
 .score_0 (score_0_x165),
 .score_1 (score_1_x165),
 .score_2 (score_2_x165),
 .score_3 (score_3_x165),
 .score_4 (score_4_x165),
 .score_5 (score_5_x165),
 .score_6 (score_6_x165),
 .score_7 (score_7_x165),
 .score_8 (score_8_x165),
 .score_9 (score_9_x165)
);
 
myram_28X28 #(
.ID(166),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x166),
.W_1(W_1_x166),
.W_2(W_2_x166),
.W_3(W_3_x166),
.W_4(W_4_x166),
.W_5(W_5_x166),
.W_6(W_6_x166),
.W_7(W_7_x166),
.W_8(W_8_x166),
.W_9(W_9_x166)
) u_28X28_x166 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x166),
 .score_0 (score_0_x166),
 .score_1 (score_1_x166),
 .score_2 (score_2_x166),
 .score_3 (score_3_x166),
 .score_4 (score_4_x166),
 .score_5 (score_5_x166),
 .score_6 (score_6_x166),
 .score_7 (score_7_x166),
 .score_8 (score_8_x166),
 .score_9 (score_9_x166)
);
 
myram_28X28 #(
.ID(167),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x167),
.W_1(W_1_x167),
.W_2(W_2_x167),
.W_3(W_3_x167),
.W_4(W_4_x167),
.W_5(W_5_x167),
.W_6(W_6_x167),
.W_7(W_7_x167),
.W_8(W_8_x167),
.W_9(W_9_x167)
) u_28X28_x167 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x167),
 .score_0 (score_0_x167),
 .score_1 (score_1_x167),
 .score_2 (score_2_x167),
 .score_3 (score_3_x167),
 .score_4 (score_4_x167),
 .score_5 (score_5_x167),
 .score_6 (score_6_x167),
 .score_7 (score_7_x167),
 .score_8 (score_8_x167),
 .score_9 (score_9_x167)
);
 
myram_28X28 #(
.ID(168),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x168),
.W_1(W_1_x168),
.W_2(W_2_x168),
.W_3(W_3_x168),
.W_4(W_4_x168),
.W_5(W_5_x168),
.W_6(W_6_x168),
.W_7(W_7_x168),
.W_8(W_8_x168),
.W_9(W_9_x168)
) u_28X28_x168 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x168),
 .score_0 (score_0_x168),
 .score_1 (score_1_x168),
 .score_2 (score_2_x168),
 .score_3 (score_3_x168),
 .score_4 (score_4_x168),
 .score_5 (score_5_x168),
 .score_6 (score_6_x168),
 .score_7 (score_7_x168),
 .score_8 (score_8_x168),
 .score_9 (score_9_x168)
);
 
myram_28X28 #(
.ID(169),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x169),
.W_1(W_1_x169),
.W_2(W_2_x169),
.W_3(W_3_x169),
.W_4(W_4_x169),
.W_5(W_5_x169),
.W_6(W_6_x169),
.W_7(W_7_x169),
.W_8(W_8_x169),
.W_9(W_9_x169)
) u_28X28_x169 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x169),
 .score_0 (score_0_x169),
 .score_1 (score_1_x169),
 .score_2 (score_2_x169),
 .score_3 (score_3_x169),
 .score_4 (score_4_x169),
 .score_5 (score_5_x169),
 .score_6 (score_6_x169),
 .score_7 (score_7_x169),
 .score_8 (score_8_x169),
 .score_9 (score_9_x169)
);
 
myram_28X28 #(
.ID(170),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x170),
.W_1(W_1_x170),
.W_2(W_2_x170),
.W_3(W_3_x170),
.W_4(W_4_x170),
.W_5(W_5_x170),
.W_6(W_6_x170),
.W_7(W_7_x170),
.W_8(W_8_x170),
.W_9(W_9_x170)
) u_28X28_x170 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x170),
 .score_0 (score_0_x170),
 .score_1 (score_1_x170),
 .score_2 (score_2_x170),
 .score_3 (score_3_x170),
 .score_4 (score_4_x170),
 .score_5 (score_5_x170),
 .score_6 (score_6_x170),
 .score_7 (score_7_x170),
 .score_8 (score_8_x170),
 .score_9 (score_9_x170)
);
 
myram_28X28 #(
.ID(171),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x171),
.W_1(W_1_x171),
.W_2(W_2_x171),
.W_3(W_3_x171),
.W_4(W_4_x171),
.W_5(W_5_x171),
.W_6(W_6_x171),
.W_7(W_7_x171),
.W_8(W_8_x171),
.W_9(W_9_x171)
) u_28X28_x171 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x171),
 .score_0 (score_0_x171),
 .score_1 (score_1_x171),
 .score_2 (score_2_x171),
 .score_3 (score_3_x171),
 .score_4 (score_4_x171),
 .score_5 (score_5_x171),
 .score_6 (score_6_x171),
 .score_7 (score_7_x171),
 .score_8 (score_8_x171),
 .score_9 (score_9_x171)
);
 
myram_28X28 #(
.ID(172),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x172),
.W_1(W_1_x172),
.W_2(W_2_x172),
.W_3(W_3_x172),
.W_4(W_4_x172),
.W_5(W_5_x172),
.W_6(W_6_x172),
.W_7(W_7_x172),
.W_8(W_8_x172),
.W_9(W_9_x172)
) u_28X28_x172 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x172),
 .score_0 (score_0_x172),
 .score_1 (score_1_x172),
 .score_2 (score_2_x172),
 .score_3 (score_3_x172),
 .score_4 (score_4_x172),
 .score_5 (score_5_x172),
 .score_6 (score_6_x172),
 .score_7 (score_7_x172),
 .score_8 (score_8_x172),
 .score_9 (score_9_x172)
);
 
myram_28X28 #(
.ID(173),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x173),
.W_1(W_1_x173),
.W_2(W_2_x173),
.W_3(W_3_x173),
.W_4(W_4_x173),
.W_5(W_5_x173),
.W_6(W_6_x173),
.W_7(W_7_x173),
.W_8(W_8_x173),
.W_9(W_9_x173)
) u_28X28_x173 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x173),
 .score_0 (score_0_x173),
 .score_1 (score_1_x173),
 .score_2 (score_2_x173),
 .score_3 (score_3_x173),
 .score_4 (score_4_x173),
 .score_5 (score_5_x173),
 .score_6 (score_6_x173),
 .score_7 (score_7_x173),
 .score_8 (score_8_x173),
 .score_9 (score_9_x173)
);
 
myram_28X28 #(
.ID(174),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x174),
.W_1(W_1_x174),
.W_2(W_2_x174),
.W_3(W_3_x174),
.W_4(W_4_x174),
.W_5(W_5_x174),
.W_6(W_6_x174),
.W_7(W_7_x174),
.W_8(W_8_x174),
.W_9(W_9_x174)
) u_28X28_x174 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x174),
 .score_0 (score_0_x174),
 .score_1 (score_1_x174),
 .score_2 (score_2_x174),
 .score_3 (score_3_x174),
 .score_4 (score_4_x174),
 .score_5 (score_5_x174),
 .score_6 (score_6_x174),
 .score_7 (score_7_x174),
 .score_8 (score_8_x174),
 .score_9 (score_9_x174)
);
 
myram_28X28 #(
.ID(175),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x175),
.W_1(W_1_x175),
.W_2(W_2_x175),
.W_3(W_3_x175),
.W_4(W_4_x175),
.W_5(W_5_x175),
.W_6(W_6_x175),
.W_7(W_7_x175),
.W_8(W_8_x175),
.W_9(W_9_x175)
) u_28X28_x175 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x175),
 .score_0 (score_0_x175),
 .score_1 (score_1_x175),
 .score_2 (score_2_x175),
 .score_3 (score_3_x175),
 .score_4 (score_4_x175),
 .score_5 (score_5_x175),
 .score_6 (score_6_x175),
 .score_7 (score_7_x175),
 .score_8 (score_8_x175),
 .score_9 (score_9_x175)
);
 
myram_28X28 #(
.ID(176),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x176),
.W_1(W_1_x176),
.W_2(W_2_x176),
.W_3(W_3_x176),
.W_4(W_4_x176),
.W_5(W_5_x176),
.W_6(W_6_x176),
.W_7(W_7_x176),
.W_8(W_8_x176),
.W_9(W_9_x176)
) u_28X28_x176 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x176),
 .score_0 (score_0_x176),
 .score_1 (score_1_x176),
 .score_2 (score_2_x176),
 .score_3 (score_3_x176),
 .score_4 (score_4_x176),
 .score_5 (score_5_x176),
 .score_6 (score_6_x176),
 .score_7 (score_7_x176),
 .score_8 (score_8_x176),
 .score_9 (score_9_x176)
);
 
myram_28X28 #(
.ID(177),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x177),
.W_1(W_1_x177),
.W_2(W_2_x177),
.W_3(W_3_x177),
.W_4(W_4_x177),
.W_5(W_5_x177),
.W_6(W_6_x177),
.W_7(W_7_x177),
.W_8(W_8_x177),
.W_9(W_9_x177)
) u_28X28_x177 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x177),
 .score_0 (score_0_x177),
 .score_1 (score_1_x177),
 .score_2 (score_2_x177),
 .score_3 (score_3_x177),
 .score_4 (score_4_x177),
 .score_5 (score_5_x177),
 .score_6 (score_6_x177),
 .score_7 (score_7_x177),
 .score_8 (score_8_x177),
 .score_9 (score_9_x177)
);
 
myram_28X28 #(
.ID(178),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x178),
.W_1(W_1_x178),
.W_2(W_2_x178),
.W_3(W_3_x178),
.W_4(W_4_x178),
.W_5(W_5_x178),
.W_6(W_6_x178),
.W_7(W_7_x178),
.W_8(W_8_x178),
.W_9(W_9_x178)
) u_28X28_x178 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x178),
 .score_0 (score_0_x178),
 .score_1 (score_1_x178),
 .score_2 (score_2_x178),
 .score_3 (score_3_x178),
 .score_4 (score_4_x178),
 .score_5 (score_5_x178),
 .score_6 (score_6_x178),
 .score_7 (score_7_x178),
 .score_8 (score_8_x178),
 .score_9 (score_9_x178)
);
 
myram_28X28 #(
.ID(179),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x179),
.W_1(W_1_x179),
.W_2(W_2_x179),
.W_3(W_3_x179),
.W_4(W_4_x179),
.W_5(W_5_x179),
.W_6(W_6_x179),
.W_7(W_7_x179),
.W_8(W_8_x179),
.W_9(W_9_x179)
) u_28X28_x179 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x179),
 .score_0 (score_0_x179),
 .score_1 (score_1_x179),
 .score_2 (score_2_x179),
 .score_3 (score_3_x179),
 .score_4 (score_4_x179),
 .score_5 (score_5_x179),
 .score_6 (score_6_x179),
 .score_7 (score_7_x179),
 .score_8 (score_8_x179),
 .score_9 (score_9_x179)
);
 
myram_28X28 #(
.ID(180),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x180),
.W_1(W_1_x180),
.W_2(W_2_x180),
.W_3(W_3_x180),
.W_4(W_4_x180),
.W_5(W_5_x180),
.W_6(W_6_x180),
.W_7(W_7_x180),
.W_8(W_8_x180),
.W_9(W_9_x180)
) u_28X28_x180 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x180),
 .score_0 (score_0_x180),
 .score_1 (score_1_x180),
 .score_2 (score_2_x180),
 .score_3 (score_3_x180),
 .score_4 (score_4_x180),
 .score_5 (score_5_x180),
 .score_6 (score_6_x180),
 .score_7 (score_7_x180),
 .score_8 (score_8_x180),
 .score_9 (score_9_x180)
);
 
myram_28X28 #(
.ID(181),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x181),
.W_1(W_1_x181),
.W_2(W_2_x181),
.W_3(W_3_x181),
.W_4(W_4_x181),
.W_5(W_5_x181),
.W_6(W_6_x181),
.W_7(W_7_x181),
.W_8(W_8_x181),
.W_9(W_9_x181)
) u_28X28_x181 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x181),
 .score_0 (score_0_x181),
 .score_1 (score_1_x181),
 .score_2 (score_2_x181),
 .score_3 (score_3_x181),
 .score_4 (score_4_x181),
 .score_5 (score_5_x181),
 .score_6 (score_6_x181),
 .score_7 (score_7_x181),
 .score_8 (score_8_x181),
 .score_9 (score_9_x181)
);
 
myram_28X28 #(
.ID(182),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x182),
.W_1(W_1_x182),
.W_2(W_2_x182),
.W_3(W_3_x182),
.W_4(W_4_x182),
.W_5(W_5_x182),
.W_6(W_6_x182),
.W_7(W_7_x182),
.W_8(W_8_x182),
.W_9(W_9_x182)
) u_28X28_x182 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x182),
 .score_0 (score_0_x182),
 .score_1 (score_1_x182),
 .score_2 (score_2_x182),
 .score_3 (score_3_x182),
 .score_4 (score_4_x182),
 .score_5 (score_5_x182),
 .score_6 (score_6_x182),
 .score_7 (score_7_x182),
 .score_8 (score_8_x182),
 .score_9 (score_9_x182)
);
 
myram_28X28 #(
.ID(183),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x183),
.W_1(W_1_x183),
.W_2(W_2_x183),
.W_3(W_3_x183),
.W_4(W_4_x183),
.W_5(W_5_x183),
.W_6(W_6_x183),
.W_7(W_7_x183),
.W_8(W_8_x183),
.W_9(W_9_x183)
) u_28X28_x183 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x183),
 .score_0 (score_0_x183),
 .score_1 (score_1_x183),
 .score_2 (score_2_x183),
 .score_3 (score_3_x183),
 .score_4 (score_4_x183),
 .score_5 (score_5_x183),
 .score_6 (score_6_x183),
 .score_7 (score_7_x183),
 .score_8 (score_8_x183),
 .score_9 (score_9_x183)
);
 
myram_28X28 #(
.ID(184),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x184),
.W_1(W_1_x184),
.W_2(W_2_x184),
.W_3(W_3_x184),
.W_4(W_4_x184),
.W_5(W_5_x184),
.W_6(W_6_x184),
.W_7(W_7_x184),
.W_8(W_8_x184),
.W_9(W_9_x184)
) u_28X28_x184 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x184),
 .score_0 (score_0_x184),
 .score_1 (score_1_x184),
 .score_2 (score_2_x184),
 .score_3 (score_3_x184),
 .score_4 (score_4_x184),
 .score_5 (score_5_x184),
 .score_6 (score_6_x184),
 .score_7 (score_7_x184),
 .score_8 (score_8_x184),
 .score_9 (score_9_x184)
);
 
myram_28X28 #(
.ID(185),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x185),
.W_1(W_1_x185),
.W_2(W_2_x185),
.W_3(W_3_x185),
.W_4(W_4_x185),
.W_5(W_5_x185),
.W_6(W_6_x185),
.W_7(W_7_x185),
.W_8(W_8_x185),
.W_9(W_9_x185)
) u_28X28_x185 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x185),
 .score_0 (score_0_x185),
 .score_1 (score_1_x185),
 .score_2 (score_2_x185),
 .score_3 (score_3_x185),
 .score_4 (score_4_x185),
 .score_5 (score_5_x185),
 .score_6 (score_6_x185),
 .score_7 (score_7_x185),
 .score_8 (score_8_x185),
 .score_9 (score_9_x185)
);
 
myram_28X28 #(
.ID(186),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x186),
.W_1(W_1_x186),
.W_2(W_2_x186),
.W_3(W_3_x186),
.W_4(W_4_x186),
.W_5(W_5_x186),
.W_6(W_6_x186),
.W_7(W_7_x186),
.W_8(W_8_x186),
.W_9(W_9_x186)
) u_28X28_x186 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x186),
 .score_0 (score_0_x186),
 .score_1 (score_1_x186),
 .score_2 (score_2_x186),
 .score_3 (score_3_x186),
 .score_4 (score_4_x186),
 .score_5 (score_5_x186),
 .score_6 (score_6_x186),
 .score_7 (score_7_x186),
 .score_8 (score_8_x186),
 .score_9 (score_9_x186)
);
 
myram_28X28 #(
.ID(187),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x187),
.W_1(W_1_x187),
.W_2(W_2_x187),
.W_3(W_3_x187),
.W_4(W_4_x187),
.W_5(W_5_x187),
.W_6(W_6_x187),
.W_7(W_7_x187),
.W_8(W_8_x187),
.W_9(W_9_x187)
) u_28X28_x187 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x187),
 .score_0 (score_0_x187),
 .score_1 (score_1_x187),
 .score_2 (score_2_x187),
 .score_3 (score_3_x187),
 .score_4 (score_4_x187),
 .score_5 (score_5_x187),
 .score_6 (score_6_x187),
 .score_7 (score_7_x187),
 .score_8 (score_8_x187),
 .score_9 (score_9_x187)
);
 
myram_28X28 #(
.ID(188),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x188),
.W_1(W_1_x188),
.W_2(W_2_x188),
.W_3(W_3_x188),
.W_4(W_4_x188),
.W_5(W_5_x188),
.W_6(W_6_x188),
.W_7(W_7_x188),
.W_8(W_8_x188),
.W_9(W_9_x188)
) u_28X28_x188 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x188),
 .score_0 (score_0_x188),
 .score_1 (score_1_x188),
 .score_2 (score_2_x188),
 .score_3 (score_3_x188),
 .score_4 (score_4_x188),
 .score_5 (score_5_x188),
 .score_6 (score_6_x188),
 .score_7 (score_7_x188),
 .score_8 (score_8_x188),
 .score_9 (score_9_x188)
);
 
myram_28X28 #(
.ID(189),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x189),
.W_1(W_1_x189),
.W_2(W_2_x189),
.W_3(W_3_x189),
.W_4(W_4_x189),
.W_5(W_5_x189),
.W_6(W_6_x189),
.W_7(W_7_x189),
.W_8(W_8_x189),
.W_9(W_9_x189)
) u_28X28_x189 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x189),
 .score_0 (score_0_x189),
 .score_1 (score_1_x189),
 .score_2 (score_2_x189),
 .score_3 (score_3_x189),
 .score_4 (score_4_x189),
 .score_5 (score_5_x189),
 .score_6 (score_6_x189),
 .score_7 (score_7_x189),
 .score_8 (score_8_x189),
 .score_9 (score_9_x189)
);
 
myram_28X28 #(
.ID(190),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x190),
.W_1(W_1_x190),
.W_2(W_2_x190),
.W_3(W_3_x190),
.W_4(W_4_x190),
.W_5(W_5_x190),
.W_6(W_6_x190),
.W_7(W_7_x190),
.W_8(W_8_x190),
.W_9(W_9_x190)
) u_28X28_x190 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x190),
 .score_0 (score_0_x190),
 .score_1 (score_1_x190),
 .score_2 (score_2_x190),
 .score_3 (score_3_x190),
 .score_4 (score_4_x190),
 .score_5 (score_5_x190),
 .score_6 (score_6_x190),
 .score_7 (score_7_x190),
 .score_8 (score_8_x190),
 .score_9 (score_9_x190)
);
 
myram_28X28 #(
.ID(191),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x191),
.W_1(W_1_x191),
.W_2(W_2_x191),
.W_3(W_3_x191),
.W_4(W_4_x191),
.W_5(W_5_x191),
.W_6(W_6_x191),
.W_7(W_7_x191),
.W_8(W_8_x191),
.W_9(W_9_x191)
) u_28X28_x191 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x191),
 .score_0 (score_0_x191),
 .score_1 (score_1_x191),
 .score_2 (score_2_x191),
 .score_3 (score_3_x191),
 .score_4 (score_4_x191),
 .score_5 (score_5_x191),
 .score_6 (score_6_x191),
 .score_7 (score_7_x191),
 .score_8 (score_8_x191),
 .score_9 (score_9_x191)
);
 
myram_28X28 #(
.ID(192),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x192),
.W_1(W_1_x192),
.W_2(W_2_x192),
.W_3(W_3_x192),
.W_4(W_4_x192),
.W_5(W_5_x192),
.W_6(W_6_x192),
.W_7(W_7_x192),
.W_8(W_8_x192),
.W_9(W_9_x192)
) u_28X28_x192 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x192),
 .score_0 (score_0_x192),
 .score_1 (score_1_x192),
 .score_2 (score_2_x192),
 .score_3 (score_3_x192),
 .score_4 (score_4_x192),
 .score_5 (score_5_x192),
 .score_6 (score_6_x192),
 .score_7 (score_7_x192),
 .score_8 (score_8_x192),
 .score_9 (score_9_x192)
);
 
myram_28X28 #(
.ID(193),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x193),
.W_1(W_1_x193),
.W_2(W_2_x193),
.W_3(W_3_x193),
.W_4(W_4_x193),
.W_5(W_5_x193),
.W_6(W_6_x193),
.W_7(W_7_x193),
.W_8(W_8_x193),
.W_9(W_9_x193)
) u_28X28_x193 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x193),
 .score_0 (score_0_x193),
 .score_1 (score_1_x193),
 .score_2 (score_2_x193),
 .score_3 (score_3_x193),
 .score_4 (score_4_x193),
 .score_5 (score_5_x193),
 .score_6 (score_6_x193),
 .score_7 (score_7_x193),
 .score_8 (score_8_x193),
 .score_9 (score_9_x193)
);
 
myram_28X28 #(
.ID(194),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x194),
.W_1(W_1_x194),
.W_2(W_2_x194),
.W_3(W_3_x194),
.W_4(W_4_x194),
.W_5(W_5_x194),
.W_6(W_6_x194),
.W_7(W_7_x194),
.W_8(W_8_x194),
.W_9(W_9_x194)
) u_28X28_x194 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x194),
 .score_0 (score_0_x194),
 .score_1 (score_1_x194),
 .score_2 (score_2_x194),
 .score_3 (score_3_x194),
 .score_4 (score_4_x194),
 .score_5 (score_5_x194),
 .score_6 (score_6_x194),
 .score_7 (score_7_x194),
 .score_8 (score_8_x194),
 .score_9 (score_9_x194)
);
 
myram_28X28 #(
.ID(195),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x195),
.W_1(W_1_x195),
.W_2(W_2_x195),
.W_3(W_3_x195),
.W_4(W_4_x195),
.W_5(W_5_x195),
.W_6(W_6_x195),
.W_7(W_7_x195),
.W_8(W_8_x195),
.W_9(W_9_x195)
) u_28X28_x195 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x195),
 .score_0 (score_0_x195),
 .score_1 (score_1_x195),
 .score_2 (score_2_x195),
 .score_3 (score_3_x195),
 .score_4 (score_4_x195),
 .score_5 (score_5_x195),
 .score_6 (score_6_x195),
 .score_7 (score_7_x195),
 .score_8 (score_8_x195),
 .score_9 (score_9_x195)
);
 
myram_28X28 #(
.ID(196),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x196),
.W_1(W_1_x196),
.W_2(W_2_x196),
.W_3(W_3_x196),
.W_4(W_4_x196),
.W_5(W_5_x196),
.W_6(W_6_x196),
.W_7(W_7_x196),
.W_8(W_8_x196),
.W_9(W_9_x196)
) u_28X28_x196 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x196),
 .score_0 (score_0_x196),
 .score_1 (score_1_x196),
 .score_2 (score_2_x196),
 .score_3 (score_3_x196),
 .score_4 (score_4_x196),
 .score_5 (score_5_x196),
 .score_6 (score_6_x196),
 .score_7 (score_7_x196),
 .score_8 (score_8_x196),
 .score_9 (score_9_x196)
);
 
myram_28X28 #(
.ID(197),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x197),
.W_1(W_1_x197),
.W_2(W_2_x197),
.W_3(W_3_x197),
.W_4(W_4_x197),
.W_5(W_5_x197),
.W_6(W_6_x197),
.W_7(W_7_x197),
.W_8(W_8_x197),
.W_9(W_9_x197)
) u_28X28_x197 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x197),
 .score_0 (score_0_x197),
 .score_1 (score_1_x197),
 .score_2 (score_2_x197),
 .score_3 (score_3_x197),
 .score_4 (score_4_x197),
 .score_5 (score_5_x197),
 .score_6 (score_6_x197),
 .score_7 (score_7_x197),
 .score_8 (score_8_x197),
 .score_9 (score_9_x197)
);
 
myram_28X28 #(
.ID(198),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x198),
.W_1(W_1_x198),
.W_2(W_2_x198),
.W_3(W_3_x198),
.W_4(W_4_x198),
.W_5(W_5_x198),
.W_6(W_6_x198),
.W_7(W_7_x198),
.W_8(W_8_x198),
.W_9(W_9_x198)
) u_28X28_x198 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x198),
 .score_0 (score_0_x198),
 .score_1 (score_1_x198),
 .score_2 (score_2_x198),
 .score_3 (score_3_x198),
 .score_4 (score_4_x198),
 .score_5 (score_5_x198),
 .score_6 (score_6_x198),
 .score_7 (score_7_x198),
 .score_8 (score_8_x198),
 .score_9 (score_9_x198)
);
 
myram_28X28 #(
.ID(199),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x199),
.W_1(W_1_x199),
.W_2(W_2_x199),
.W_3(W_3_x199),
.W_4(W_4_x199),
.W_5(W_5_x199),
.W_6(W_6_x199),
.W_7(W_7_x199),
.W_8(W_8_x199),
.W_9(W_9_x199)
) u_28X28_x199 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x199),
 .score_0 (score_0_x199),
 .score_1 (score_1_x199),
 .score_2 (score_2_x199),
 .score_3 (score_3_x199),
 .score_4 (score_4_x199),
 .score_5 (score_5_x199),
 .score_6 (score_6_x199),
 .score_7 (score_7_x199),
 .score_8 (score_8_x199),
 .score_9 (score_9_x199)
);
 
myram_28X28 #(
.ID(200),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x200),
.W_1(W_1_x200),
.W_2(W_2_x200),
.W_3(W_3_x200),
.W_4(W_4_x200),
.W_5(W_5_x200),
.W_6(W_6_x200),
.W_7(W_7_x200),
.W_8(W_8_x200),
.W_9(W_9_x200)
) u_28X28_x200 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x200),
 .score_0 (score_0_x200),
 .score_1 (score_1_x200),
 .score_2 (score_2_x200),
 .score_3 (score_3_x200),
 .score_4 (score_4_x200),
 .score_5 (score_5_x200),
 .score_6 (score_6_x200),
 .score_7 (score_7_x200),
 .score_8 (score_8_x200),
 .score_9 (score_9_x200)
);
 
myram_28X28 #(
.ID(201),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x201),
.W_1(W_1_x201),
.W_2(W_2_x201),
.W_3(W_3_x201),
.W_4(W_4_x201),
.W_5(W_5_x201),
.W_6(W_6_x201),
.W_7(W_7_x201),
.W_8(W_8_x201),
.W_9(W_9_x201)
) u_28X28_x201 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x201),
 .score_0 (score_0_x201),
 .score_1 (score_1_x201),
 .score_2 (score_2_x201),
 .score_3 (score_3_x201),
 .score_4 (score_4_x201),
 .score_5 (score_5_x201),
 .score_6 (score_6_x201),
 .score_7 (score_7_x201),
 .score_8 (score_8_x201),
 .score_9 (score_9_x201)
);
 
myram_28X28 #(
.ID(202),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x202),
.W_1(W_1_x202),
.W_2(W_2_x202),
.W_3(W_3_x202),
.W_4(W_4_x202),
.W_5(W_5_x202),
.W_6(W_6_x202),
.W_7(W_7_x202),
.W_8(W_8_x202),
.W_9(W_9_x202)
) u_28X28_x202 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x202),
 .score_0 (score_0_x202),
 .score_1 (score_1_x202),
 .score_2 (score_2_x202),
 .score_3 (score_3_x202),
 .score_4 (score_4_x202),
 .score_5 (score_5_x202),
 .score_6 (score_6_x202),
 .score_7 (score_7_x202),
 .score_8 (score_8_x202),
 .score_9 (score_9_x202)
);
 
myram_28X28 #(
.ID(203),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x203),
.W_1(W_1_x203),
.W_2(W_2_x203),
.W_3(W_3_x203),
.W_4(W_4_x203),
.W_5(W_5_x203),
.W_6(W_6_x203),
.W_7(W_7_x203),
.W_8(W_8_x203),
.W_9(W_9_x203)
) u_28X28_x203 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x203),
 .score_0 (score_0_x203),
 .score_1 (score_1_x203),
 .score_2 (score_2_x203),
 .score_3 (score_3_x203),
 .score_4 (score_4_x203),
 .score_5 (score_5_x203),
 .score_6 (score_6_x203),
 .score_7 (score_7_x203),
 .score_8 (score_8_x203),
 .score_9 (score_9_x203)
);
 
myram_28X28 #(
.ID(204),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x204),
.W_1(W_1_x204),
.W_2(W_2_x204),
.W_3(W_3_x204),
.W_4(W_4_x204),
.W_5(W_5_x204),
.W_6(W_6_x204),
.W_7(W_7_x204),
.W_8(W_8_x204),
.W_9(W_9_x204)
) u_28X28_x204 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x204),
 .score_0 (score_0_x204),
 .score_1 (score_1_x204),
 .score_2 (score_2_x204),
 .score_3 (score_3_x204),
 .score_4 (score_4_x204),
 .score_5 (score_5_x204),
 .score_6 (score_6_x204),
 .score_7 (score_7_x204),
 .score_8 (score_8_x204),
 .score_9 (score_9_x204)
);
 
myram_28X28 #(
.ID(205),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x205),
.W_1(W_1_x205),
.W_2(W_2_x205),
.W_3(W_3_x205),
.W_4(W_4_x205),
.W_5(W_5_x205),
.W_6(W_6_x205),
.W_7(W_7_x205),
.W_8(W_8_x205),
.W_9(W_9_x205)
) u_28X28_x205 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x205),
 .score_0 (score_0_x205),
 .score_1 (score_1_x205),
 .score_2 (score_2_x205),
 .score_3 (score_3_x205),
 .score_4 (score_4_x205),
 .score_5 (score_5_x205),
 .score_6 (score_6_x205),
 .score_7 (score_7_x205),
 .score_8 (score_8_x205),
 .score_9 (score_9_x205)
);
 
myram_28X28 #(
.ID(206),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x206),
.W_1(W_1_x206),
.W_2(W_2_x206),
.W_3(W_3_x206),
.W_4(W_4_x206),
.W_5(W_5_x206),
.W_6(W_6_x206),
.W_7(W_7_x206),
.W_8(W_8_x206),
.W_9(W_9_x206)
) u_28X28_x206 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x206),
 .score_0 (score_0_x206),
 .score_1 (score_1_x206),
 .score_2 (score_2_x206),
 .score_3 (score_3_x206),
 .score_4 (score_4_x206),
 .score_5 (score_5_x206),
 .score_6 (score_6_x206),
 .score_7 (score_7_x206),
 .score_8 (score_8_x206),
 .score_9 (score_9_x206)
);
 
myram_28X28 #(
.ID(207),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x207),
.W_1(W_1_x207),
.W_2(W_2_x207),
.W_3(W_3_x207),
.W_4(W_4_x207),
.W_5(W_5_x207),
.W_6(W_6_x207),
.W_7(W_7_x207),
.W_8(W_8_x207),
.W_9(W_9_x207)
) u_28X28_x207 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x207),
 .score_0 (score_0_x207),
 .score_1 (score_1_x207),
 .score_2 (score_2_x207),
 .score_3 (score_3_x207),
 .score_4 (score_4_x207),
 .score_5 (score_5_x207),
 .score_6 (score_6_x207),
 .score_7 (score_7_x207),
 .score_8 (score_8_x207),
 .score_9 (score_9_x207)
);
 
myram_28X28 #(
.ID(208),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x208),
.W_1(W_1_x208),
.W_2(W_2_x208),
.W_3(W_3_x208),
.W_4(W_4_x208),
.W_5(W_5_x208),
.W_6(W_6_x208),
.W_7(W_7_x208),
.W_8(W_8_x208),
.W_9(W_9_x208)
) u_28X28_x208 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x208),
 .score_0 (score_0_x208),
 .score_1 (score_1_x208),
 .score_2 (score_2_x208),
 .score_3 (score_3_x208),
 .score_4 (score_4_x208),
 .score_5 (score_5_x208),
 .score_6 (score_6_x208),
 .score_7 (score_7_x208),
 .score_8 (score_8_x208),
 .score_9 (score_9_x208)
);
 
myram_28X28 #(
.ID(209),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x209),
.W_1(W_1_x209),
.W_2(W_2_x209),
.W_3(W_3_x209),
.W_4(W_4_x209),
.W_5(W_5_x209),
.W_6(W_6_x209),
.W_7(W_7_x209),
.W_8(W_8_x209),
.W_9(W_9_x209)
) u_28X28_x209 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x209),
 .score_0 (score_0_x209),
 .score_1 (score_1_x209),
 .score_2 (score_2_x209),
 .score_3 (score_3_x209),
 .score_4 (score_4_x209),
 .score_5 (score_5_x209),
 .score_6 (score_6_x209),
 .score_7 (score_7_x209),
 .score_8 (score_8_x209),
 .score_9 (score_9_x209)
);
 
myram_28X28 #(
.ID(210),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x210),
.W_1(W_1_x210),
.W_2(W_2_x210),
.W_3(W_3_x210),
.W_4(W_4_x210),
.W_5(W_5_x210),
.W_6(W_6_x210),
.W_7(W_7_x210),
.W_8(W_8_x210),
.W_9(W_9_x210)
) u_28X28_x210 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x210),
 .score_0 (score_0_x210),
 .score_1 (score_1_x210),
 .score_2 (score_2_x210),
 .score_3 (score_3_x210),
 .score_4 (score_4_x210),
 .score_5 (score_5_x210),
 .score_6 (score_6_x210),
 .score_7 (score_7_x210),
 .score_8 (score_8_x210),
 .score_9 (score_9_x210)
);
 
myram_28X28 #(
.ID(211),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x211),
.W_1(W_1_x211),
.W_2(W_2_x211),
.W_3(W_3_x211),
.W_4(W_4_x211),
.W_5(W_5_x211),
.W_6(W_6_x211),
.W_7(W_7_x211),
.W_8(W_8_x211),
.W_9(W_9_x211)
) u_28X28_x211 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x211),
 .score_0 (score_0_x211),
 .score_1 (score_1_x211),
 .score_2 (score_2_x211),
 .score_3 (score_3_x211),
 .score_4 (score_4_x211),
 .score_5 (score_5_x211),
 .score_6 (score_6_x211),
 .score_7 (score_7_x211),
 .score_8 (score_8_x211),
 .score_9 (score_9_x211)
);
 
myram_28X28 #(
.ID(212),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x212),
.W_1(W_1_x212),
.W_2(W_2_x212),
.W_3(W_3_x212),
.W_4(W_4_x212),
.W_5(W_5_x212),
.W_6(W_6_x212),
.W_7(W_7_x212),
.W_8(W_8_x212),
.W_9(W_9_x212)
) u_28X28_x212 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x212),
 .score_0 (score_0_x212),
 .score_1 (score_1_x212),
 .score_2 (score_2_x212),
 .score_3 (score_3_x212),
 .score_4 (score_4_x212),
 .score_5 (score_5_x212),
 .score_6 (score_6_x212),
 .score_7 (score_7_x212),
 .score_8 (score_8_x212),
 .score_9 (score_9_x212)
);
 
myram_28X28 #(
.ID(213),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x213),
.W_1(W_1_x213),
.W_2(W_2_x213),
.W_3(W_3_x213),
.W_4(W_4_x213),
.W_5(W_5_x213),
.W_6(W_6_x213),
.W_7(W_7_x213),
.W_8(W_8_x213),
.W_9(W_9_x213)
) u_28X28_x213 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x213),
 .score_0 (score_0_x213),
 .score_1 (score_1_x213),
 .score_2 (score_2_x213),
 .score_3 (score_3_x213),
 .score_4 (score_4_x213),
 .score_5 (score_5_x213),
 .score_6 (score_6_x213),
 .score_7 (score_7_x213),
 .score_8 (score_8_x213),
 .score_9 (score_9_x213)
);
 
myram_28X28 #(
.ID(214),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x214),
.W_1(W_1_x214),
.W_2(W_2_x214),
.W_3(W_3_x214),
.W_4(W_4_x214),
.W_5(W_5_x214),
.W_6(W_6_x214),
.W_7(W_7_x214),
.W_8(W_8_x214),
.W_9(W_9_x214)
) u_28X28_x214 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x214),
 .score_0 (score_0_x214),
 .score_1 (score_1_x214),
 .score_2 (score_2_x214),
 .score_3 (score_3_x214),
 .score_4 (score_4_x214),
 .score_5 (score_5_x214),
 .score_6 (score_6_x214),
 .score_7 (score_7_x214),
 .score_8 (score_8_x214),
 .score_9 (score_9_x214)
);
 
myram_28X28 #(
.ID(215),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x215),
.W_1(W_1_x215),
.W_2(W_2_x215),
.W_3(W_3_x215),
.W_4(W_4_x215),
.W_5(W_5_x215),
.W_6(W_6_x215),
.W_7(W_7_x215),
.W_8(W_8_x215),
.W_9(W_9_x215)
) u_28X28_x215 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x215),
 .score_0 (score_0_x215),
 .score_1 (score_1_x215),
 .score_2 (score_2_x215),
 .score_3 (score_3_x215),
 .score_4 (score_4_x215),
 .score_5 (score_5_x215),
 .score_6 (score_6_x215),
 .score_7 (score_7_x215),
 .score_8 (score_8_x215),
 .score_9 (score_9_x215)
);
 
myram_28X28 #(
.ID(216),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x216),
.W_1(W_1_x216),
.W_2(W_2_x216),
.W_3(W_3_x216),
.W_4(W_4_x216),
.W_5(W_5_x216),
.W_6(W_6_x216),
.W_7(W_7_x216),
.W_8(W_8_x216),
.W_9(W_9_x216)
) u_28X28_x216 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x216),
 .score_0 (score_0_x216),
 .score_1 (score_1_x216),
 .score_2 (score_2_x216),
 .score_3 (score_3_x216),
 .score_4 (score_4_x216),
 .score_5 (score_5_x216),
 .score_6 (score_6_x216),
 .score_7 (score_7_x216),
 .score_8 (score_8_x216),
 .score_9 (score_9_x216)
);
 
myram_28X28 #(
.ID(217),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x217),
.W_1(W_1_x217),
.W_2(W_2_x217),
.W_3(W_3_x217),
.W_4(W_4_x217),
.W_5(W_5_x217),
.W_6(W_6_x217),
.W_7(W_7_x217),
.W_8(W_8_x217),
.W_9(W_9_x217)
) u_28X28_x217 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x217),
 .score_0 (score_0_x217),
 .score_1 (score_1_x217),
 .score_2 (score_2_x217),
 .score_3 (score_3_x217),
 .score_4 (score_4_x217),
 .score_5 (score_5_x217),
 .score_6 (score_6_x217),
 .score_7 (score_7_x217),
 .score_8 (score_8_x217),
 .score_9 (score_9_x217)
);
 
myram_28X28 #(
.ID(218),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x218),
.W_1(W_1_x218),
.W_2(W_2_x218),
.W_3(W_3_x218),
.W_4(W_4_x218),
.W_5(W_5_x218),
.W_6(W_6_x218),
.W_7(W_7_x218),
.W_8(W_8_x218),
.W_9(W_9_x218)
) u_28X28_x218 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x218),
 .score_0 (score_0_x218),
 .score_1 (score_1_x218),
 .score_2 (score_2_x218),
 .score_3 (score_3_x218),
 .score_4 (score_4_x218),
 .score_5 (score_5_x218),
 .score_6 (score_6_x218),
 .score_7 (score_7_x218),
 .score_8 (score_8_x218),
 .score_9 (score_9_x218)
);
 
myram_28X28 #(
.ID(219),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x219),
.W_1(W_1_x219),
.W_2(W_2_x219),
.W_3(W_3_x219),
.W_4(W_4_x219),
.W_5(W_5_x219),
.W_6(W_6_x219),
.W_7(W_7_x219),
.W_8(W_8_x219),
.W_9(W_9_x219)
) u_28X28_x219 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x219),
 .score_0 (score_0_x219),
 .score_1 (score_1_x219),
 .score_2 (score_2_x219),
 .score_3 (score_3_x219),
 .score_4 (score_4_x219),
 .score_5 (score_5_x219),
 .score_6 (score_6_x219),
 .score_7 (score_7_x219),
 .score_8 (score_8_x219),
 .score_9 (score_9_x219)
);
 
myram_28X28 #(
.ID(220),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x220),
.W_1(W_1_x220),
.W_2(W_2_x220),
.W_3(W_3_x220),
.W_4(W_4_x220),
.W_5(W_5_x220),
.W_6(W_6_x220),
.W_7(W_7_x220),
.W_8(W_8_x220),
.W_9(W_9_x220)
) u_28X28_x220 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x220),
 .score_0 (score_0_x220),
 .score_1 (score_1_x220),
 .score_2 (score_2_x220),
 .score_3 (score_3_x220),
 .score_4 (score_4_x220),
 .score_5 (score_5_x220),
 .score_6 (score_6_x220),
 .score_7 (score_7_x220),
 .score_8 (score_8_x220),
 .score_9 (score_9_x220)
);
 
myram_28X28 #(
.ID(221),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x221),
.W_1(W_1_x221),
.W_2(W_2_x221),
.W_3(W_3_x221),
.W_4(W_4_x221),
.W_5(W_5_x221),
.W_6(W_6_x221),
.W_7(W_7_x221),
.W_8(W_8_x221),
.W_9(W_9_x221)
) u_28X28_x221 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x221),
 .score_0 (score_0_x221),
 .score_1 (score_1_x221),
 .score_2 (score_2_x221),
 .score_3 (score_3_x221),
 .score_4 (score_4_x221),
 .score_5 (score_5_x221),
 .score_6 (score_6_x221),
 .score_7 (score_7_x221),
 .score_8 (score_8_x221),
 .score_9 (score_9_x221)
);
 
myram_28X28 #(
.ID(222),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x222),
.W_1(W_1_x222),
.W_2(W_2_x222),
.W_3(W_3_x222),
.W_4(W_4_x222),
.W_5(W_5_x222),
.W_6(W_6_x222),
.W_7(W_7_x222),
.W_8(W_8_x222),
.W_9(W_9_x222)
) u_28X28_x222 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x222),
 .score_0 (score_0_x222),
 .score_1 (score_1_x222),
 .score_2 (score_2_x222),
 .score_3 (score_3_x222),
 .score_4 (score_4_x222),
 .score_5 (score_5_x222),
 .score_6 (score_6_x222),
 .score_7 (score_7_x222),
 .score_8 (score_8_x222),
 .score_9 (score_9_x222)
);
 
myram_28X28 #(
.ID(223),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x223),
.W_1(W_1_x223),
.W_2(W_2_x223),
.W_3(W_3_x223),
.W_4(W_4_x223),
.W_5(W_5_x223),
.W_6(W_6_x223),
.W_7(W_7_x223),
.W_8(W_8_x223),
.W_9(W_9_x223)
) u_28X28_x223 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x223),
 .score_0 (score_0_x223),
 .score_1 (score_1_x223),
 .score_2 (score_2_x223),
 .score_3 (score_3_x223),
 .score_4 (score_4_x223),
 .score_5 (score_5_x223),
 .score_6 (score_6_x223),
 .score_7 (score_7_x223),
 .score_8 (score_8_x223),
 .score_9 (score_9_x223)
);
 
myram_28X28 #(
.ID(224),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x224),
.W_1(W_1_x224),
.W_2(W_2_x224),
.W_3(W_3_x224),
.W_4(W_4_x224),
.W_5(W_5_x224),
.W_6(W_6_x224),
.W_7(W_7_x224),
.W_8(W_8_x224),
.W_9(W_9_x224)
) u_28X28_x224 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x224),
 .score_0 (score_0_x224),
 .score_1 (score_1_x224),
 .score_2 (score_2_x224),
 .score_3 (score_3_x224),
 .score_4 (score_4_x224),
 .score_5 (score_5_x224),
 .score_6 (score_6_x224),
 .score_7 (score_7_x224),
 .score_8 (score_8_x224),
 .score_9 (score_9_x224)
);
 
myram_28X28 #(
.ID(225),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x225),
.W_1(W_1_x225),
.W_2(W_2_x225),
.W_3(W_3_x225),
.W_4(W_4_x225),
.W_5(W_5_x225),
.W_6(W_6_x225),
.W_7(W_7_x225),
.W_8(W_8_x225),
.W_9(W_9_x225)
) u_28X28_x225 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x225),
 .score_0 (score_0_x225),
 .score_1 (score_1_x225),
 .score_2 (score_2_x225),
 .score_3 (score_3_x225),
 .score_4 (score_4_x225),
 .score_5 (score_5_x225),
 .score_6 (score_6_x225),
 .score_7 (score_7_x225),
 .score_8 (score_8_x225),
 .score_9 (score_9_x225)
);
 
myram_28X28 #(
.ID(226),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x226),
.W_1(W_1_x226),
.W_2(W_2_x226),
.W_3(W_3_x226),
.W_4(W_4_x226),
.W_5(W_5_x226),
.W_6(W_6_x226),
.W_7(W_7_x226),
.W_8(W_8_x226),
.W_9(W_9_x226)
) u_28X28_x226 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x226),
 .score_0 (score_0_x226),
 .score_1 (score_1_x226),
 .score_2 (score_2_x226),
 .score_3 (score_3_x226),
 .score_4 (score_4_x226),
 .score_5 (score_5_x226),
 .score_6 (score_6_x226),
 .score_7 (score_7_x226),
 .score_8 (score_8_x226),
 .score_9 (score_9_x226)
);
 
myram_28X28 #(
.ID(227),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x227),
.W_1(W_1_x227),
.W_2(W_2_x227),
.W_3(W_3_x227),
.W_4(W_4_x227),
.W_5(W_5_x227),
.W_6(W_6_x227),
.W_7(W_7_x227),
.W_8(W_8_x227),
.W_9(W_9_x227)
) u_28X28_x227 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x227),
 .score_0 (score_0_x227),
 .score_1 (score_1_x227),
 .score_2 (score_2_x227),
 .score_3 (score_3_x227),
 .score_4 (score_4_x227),
 .score_5 (score_5_x227),
 .score_6 (score_6_x227),
 .score_7 (score_7_x227),
 .score_8 (score_8_x227),
 .score_9 (score_9_x227)
);
 
myram_28X28 #(
.ID(228),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x228),
.W_1(W_1_x228),
.W_2(W_2_x228),
.W_3(W_3_x228),
.W_4(W_4_x228),
.W_5(W_5_x228),
.W_6(W_6_x228),
.W_7(W_7_x228),
.W_8(W_8_x228),
.W_9(W_9_x228)
) u_28X28_x228 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x228),
 .score_0 (score_0_x228),
 .score_1 (score_1_x228),
 .score_2 (score_2_x228),
 .score_3 (score_3_x228),
 .score_4 (score_4_x228),
 .score_5 (score_5_x228),
 .score_6 (score_6_x228),
 .score_7 (score_7_x228),
 .score_8 (score_8_x228),
 .score_9 (score_9_x228)
);
 
myram_28X28 #(
.ID(229),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x229),
.W_1(W_1_x229),
.W_2(W_2_x229),
.W_3(W_3_x229),
.W_4(W_4_x229),
.W_5(W_5_x229),
.W_6(W_6_x229),
.W_7(W_7_x229),
.W_8(W_8_x229),
.W_9(W_9_x229)
) u_28X28_x229 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x229),
 .score_0 (score_0_x229),
 .score_1 (score_1_x229),
 .score_2 (score_2_x229),
 .score_3 (score_3_x229),
 .score_4 (score_4_x229),
 .score_5 (score_5_x229),
 .score_6 (score_6_x229),
 .score_7 (score_7_x229),
 .score_8 (score_8_x229),
 .score_9 (score_9_x229)
);
 
myram_28X28 #(
.ID(230),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x230),
.W_1(W_1_x230),
.W_2(W_2_x230),
.W_3(W_3_x230),
.W_4(W_4_x230),
.W_5(W_5_x230),
.W_6(W_6_x230),
.W_7(W_7_x230),
.W_8(W_8_x230),
.W_9(W_9_x230)
) u_28X28_x230 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x230),
 .score_0 (score_0_x230),
 .score_1 (score_1_x230),
 .score_2 (score_2_x230),
 .score_3 (score_3_x230),
 .score_4 (score_4_x230),
 .score_5 (score_5_x230),
 .score_6 (score_6_x230),
 .score_7 (score_7_x230),
 .score_8 (score_8_x230),
 .score_9 (score_9_x230)
);
 
myram_28X28 #(
.ID(231),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x231),
.W_1(W_1_x231),
.W_2(W_2_x231),
.W_3(W_3_x231),
.W_4(W_4_x231),
.W_5(W_5_x231),
.W_6(W_6_x231),
.W_7(W_7_x231),
.W_8(W_8_x231),
.W_9(W_9_x231)
) u_28X28_x231 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x231),
 .score_0 (score_0_x231),
 .score_1 (score_1_x231),
 .score_2 (score_2_x231),
 .score_3 (score_3_x231),
 .score_4 (score_4_x231),
 .score_5 (score_5_x231),
 .score_6 (score_6_x231),
 .score_7 (score_7_x231),
 .score_8 (score_8_x231),
 .score_9 (score_9_x231)
);
 
myram_28X28 #(
.ID(232),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x232),
.W_1(W_1_x232),
.W_2(W_2_x232),
.W_3(W_3_x232),
.W_4(W_4_x232),
.W_5(W_5_x232),
.W_6(W_6_x232),
.W_7(W_7_x232),
.W_8(W_8_x232),
.W_9(W_9_x232)
) u_28X28_x232 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x232),
 .score_0 (score_0_x232),
 .score_1 (score_1_x232),
 .score_2 (score_2_x232),
 .score_3 (score_3_x232),
 .score_4 (score_4_x232),
 .score_5 (score_5_x232),
 .score_6 (score_6_x232),
 .score_7 (score_7_x232),
 .score_8 (score_8_x232),
 .score_9 (score_9_x232)
);
 
myram_28X28 #(
.ID(233),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x233),
.W_1(W_1_x233),
.W_2(W_2_x233),
.W_3(W_3_x233),
.W_4(W_4_x233),
.W_5(W_5_x233),
.W_6(W_6_x233),
.W_7(W_7_x233),
.W_8(W_8_x233),
.W_9(W_9_x233)
) u_28X28_x233 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x233),
 .score_0 (score_0_x233),
 .score_1 (score_1_x233),
 .score_2 (score_2_x233),
 .score_3 (score_3_x233),
 .score_4 (score_4_x233),
 .score_5 (score_5_x233),
 .score_6 (score_6_x233),
 .score_7 (score_7_x233),
 .score_8 (score_8_x233),
 .score_9 (score_9_x233)
);
 
myram_28X28 #(
.ID(234),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x234),
.W_1(W_1_x234),
.W_2(W_2_x234),
.W_3(W_3_x234),
.W_4(W_4_x234),
.W_5(W_5_x234),
.W_6(W_6_x234),
.W_7(W_7_x234),
.W_8(W_8_x234),
.W_9(W_9_x234)
) u_28X28_x234 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x234),
 .score_0 (score_0_x234),
 .score_1 (score_1_x234),
 .score_2 (score_2_x234),
 .score_3 (score_3_x234),
 .score_4 (score_4_x234),
 .score_5 (score_5_x234),
 .score_6 (score_6_x234),
 .score_7 (score_7_x234),
 .score_8 (score_8_x234),
 .score_9 (score_9_x234)
);
 
myram_28X28 #(
.ID(235),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x235),
.W_1(W_1_x235),
.W_2(W_2_x235),
.W_3(W_3_x235),
.W_4(W_4_x235),
.W_5(W_5_x235),
.W_6(W_6_x235),
.W_7(W_7_x235),
.W_8(W_8_x235),
.W_9(W_9_x235)
) u_28X28_x235 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x235),
 .score_0 (score_0_x235),
 .score_1 (score_1_x235),
 .score_2 (score_2_x235),
 .score_3 (score_3_x235),
 .score_4 (score_4_x235),
 .score_5 (score_5_x235),
 .score_6 (score_6_x235),
 .score_7 (score_7_x235),
 .score_8 (score_8_x235),
 .score_9 (score_9_x235)
);
 
myram_28X28 #(
.ID(236),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x236),
.W_1(W_1_x236),
.W_2(W_2_x236),
.W_3(W_3_x236),
.W_4(W_4_x236),
.W_5(W_5_x236),
.W_6(W_6_x236),
.W_7(W_7_x236),
.W_8(W_8_x236),
.W_9(W_9_x236)
) u_28X28_x236 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x236),
 .score_0 (score_0_x236),
 .score_1 (score_1_x236),
 .score_2 (score_2_x236),
 .score_3 (score_3_x236),
 .score_4 (score_4_x236),
 .score_5 (score_5_x236),
 .score_6 (score_6_x236),
 .score_7 (score_7_x236),
 .score_8 (score_8_x236),
 .score_9 (score_9_x236)
);
 
myram_28X28 #(
.ID(237),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x237),
.W_1(W_1_x237),
.W_2(W_2_x237),
.W_3(W_3_x237),
.W_4(W_4_x237),
.W_5(W_5_x237),
.W_6(W_6_x237),
.W_7(W_7_x237),
.W_8(W_8_x237),
.W_9(W_9_x237)
) u_28X28_x237 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x237),
 .score_0 (score_0_x237),
 .score_1 (score_1_x237),
 .score_2 (score_2_x237),
 .score_3 (score_3_x237),
 .score_4 (score_4_x237),
 .score_5 (score_5_x237),
 .score_6 (score_6_x237),
 .score_7 (score_7_x237),
 .score_8 (score_8_x237),
 .score_9 (score_9_x237)
);
 
myram_28X28 #(
.ID(238),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x238),
.W_1(W_1_x238),
.W_2(W_2_x238),
.W_3(W_3_x238),
.W_4(W_4_x238),
.W_5(W_5_x238),
.W_6(W_6_x238),
.W_7(W_7_x238),
.W_8(W_8_x238),
.W_9(W_9_x238)
) u_28X28_x238 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x238),
 .score_0 (score_0_x238),
 .score_1 (score_1_x238),
 .score_2 (score_2_x238),
 .score_3 (score_3_x238),
 .score_4 (score_4_x238),
 .score_5 (score_5_x238),
 .score_6 (score_6_x238),
 .score_7 (score_7_x238),
 .score_8 (score_8_x238),
 .score_9 (score_9_x238)
);
 
myram_28X28 #(
.ID(239),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x239),
.W_1(W_1_x239),
.W_2(W_2_x239),
.W_3(W_3_x239),
.W_4(W_4_x239),
.W_5(W_5_x239),
.W_6(W_6_x239),
.W_7(W_7_x239),
.W_8(W_8_x239),
.W_9(W_9_x239)
) u_28X28_x239 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x239),
 .score_0 (score_0_x239),
 .score_1 (score_1_x239),
 .score_2 (score_2_x239),
 .score_3 (score_3_x239),
 .score_4 (score_4_x239),
 .score_5 (score_5_x239),
 .score_6 (score_6_x239),
 .score_7 (score_7_x239),
 .score_8 (score_8_x239),
 .score_9 (score_9_x239)
);
 
myram_28X28 #(
.ID(240),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x240),
.W_1(W_1_x240),
.W_2(W_2_x240),
.W_3(W_3_x240),
.W_4(W_4_x240),
.W_5(W_5_x240),
.W_6(W_6_x240),
.W_7(W_7_x240),
.W_8(W_8_x240),
.W_9(W_9_x240)
) u_28X28_x240 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x240),
 .score_0 (score_0_x240),
 .score_1 (score_1_x240),
 .score_2 (score_2_x240),
 .score_3 (score_3_x240),
 .score_4 (score_4_x240),
 .score_5 (score_5_x240),
 .score_6 (score_6_x240),
 .score_7 (score_7_x240),
 .score_8 (score_8_x240),
 .score_9 (score_9_x240)
);
 
myram_28X28 #(
.ID(241),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x241),
.W_1(W_1_x241),
.W_2(W_2_x241),
.W_3(W_3_x241),
.W_4(W_4_x241),
.W_5(W_5_x241),
.W_6(W_6_x241),
.W_7(W_7_x241),
.W_8(W_8_x241),
.W_9(W_9_x241)
) u_28X28_x241 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x241),
 .score_0 (score_0_x241),
 .score_1 (score_1_x241),
 .score_2 (score_2_x241),
 .score_3 (score_3_x241),
 .score_4 (score_4_x241),
 .score_5 (score_5_x241),
 .score_6 (score_6_x241),
 .score_7 (score_7_x241),
 .score_8 (score_8_x241),
 .score_9 (score_9_x241)
);
 
myram_28X28 #(
.ID(242),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x242),
.W_1(W_1_x242),
.W_2(W_2_x242),
.W_3(W_3_x242),
.W_4(W_4_x242),
.W_5(W_5_x242),
.W_6(W_6_x242),
.W_7(W_7_x242),
.W_8(W_8_x242),
.W_9(W_9_x242)
) u_28X28_x242 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x242),
 .score_0 (score_0_x242),
 .score_1 (score_1_x242),
 .score_2 (score_2_x242),
 .score_3 (score_3_x242),
 .score_4 (score_4_x242),
 .score_5 (score_5_x242),
 .score_6 (score_6_x242),
 .score_7 (score_7_x242),
 .score_8 (score_8_x242),
 .score_9 (score_9_x242)
);
 
myram_28X28 #(
.ID(243),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x243),
.W_1(W_1_x243),
.W_2(W_2_x243),
.W_3(W_3_x243),
.W_4(W_4_x243),
.W_5(W_5_x243),
.W_6(W_6_x243),
.W_7(W_7_x243),
.W_8(W_8_x243),
.W_9(W_9_x243)
) u_28X28_x243 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x243),
 .score_0 (score_0_x243),
 .score_1 (score_1_x243),
 .score_2 (score_2_x243),
 .score_3 (score_3_x243),
 .score_4 (score_4_x243),
 .score_5 (score_5_x243),
 .score_6 (score_6_x243),
 .score_7 (score_7_x243),
 .score_8 (score_8_x243),
 .score_9 (score_9_x243)
);
 
myram_28X28 #(
.ID(244),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x244),
.W_1(W_1_x244),
.W_2(W_2_x244),
.W_3(W_3_x244),
.W_4(W_4_x244),
.W_5(W_5_x244),
.W_6(W_6_x244),
.W_7(W_7_x244),
.W_8(W_8_x244),
.W_9(W_9_x244)
) u_28X28_x244 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x244),
 .score_0 (score_0_x244),
 .score_1 (score_1_x244),
 .score_2 (score_2_x244),
 .score_3 (score_3_x244),
 .score_4 (score_4_x244),
 .score_5 (score_5_x244),
 .score_6 (score_6_x244),
 .score_7 (score_7_x244),
 .score_8 (score_8_x244),
 .score_9 (score_9_x244)
);
 
myram_28X28 #(
.ID(245),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x245),
.W_1(W_1_x245),
.W_2(W_2_x245),
.W_3(W_3_x245),
.W_4(W_4_x245),
.W_5(W_5_x245),
.W_6(W_6_x245),
.W_7(W_7_x245),
.W_8(W_8_x245),
.W_9(W_9_x245)
) u_28X28_x245 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x245),
 .score_0 (score_0_x245),
 .score_1 (score_1_x245),
 .score_2 (score_2_x245),
 .score_3 (score_3_x245),
 .score_4 (score_4_x245),
 .score_5 (score_5_x245),
 .score_6 (score_6_x245),
 .score_7 (score_7_x245),
 .score_8 (score_8_x245),
 .score_9 (score_9_x245)
);
 
myram_28X28 #(
.ID(246),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x246),
.W_1(W_1_x246),
.W_2(W_2_x246),
.W_3(W_3_x246),
.W_4(W_4_x246),
.W_5(W_5_x246),
.W_6(W_6_x246),
.W_7(W_7_x246),
.W_8(W_8_x246),
.W_9(W_9_x246)
) u_28X28_x246 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x246),
 .score_0 (score_0_x246),
 .score_1 (score_1_x246),
 .score_2 (score_2_x246),
 .score_3 (score_3_x246),
 .score_4 (score_4_x246),
 .score_5 (score_5_x246),
 .score_6 (score_6_x246),
 .score_7 (score_7_x246),
 .score_8 (score_8_x246),
 .score_9 (score_9_x246)
);
 
myram_28X28 #(
.ID(247),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x247),
.W_1(W_1_x247),
.W_2(W_2_x247),
.W_3(W_3_x247),
.W_4(W_4_x247),
.W_5(W_5_x247),
.W_6(W_6_x247),
.W_7(W_7_x247),
.W_8(W_8_x247),
.W_9(W_9_x247)
) u_28X28_x247 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x247),
 .score_0 (score_0_x247),
 .score_1 (score_1_x247),
 .score_2 (score_2_x247),
 .score_3 (score_3_x247),
 .score_4 (score_4_x247),
 .score_5 (score_5_x247),
 .score_6 (score_6_x247),
 .score_7 (score_7_x247),
 .score_8 (score_8_x247),
 .score_9 (score_9_x247)
);
 
myram_28X28 #(
.ID(248),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x248),
.W_1(W_1_x248),
.W_2(W_2_x248),
.W_3(W_3_x248),
.W_4(W_4_x248),
.W_5(W_5_x248),
.W_6(W_6_x248),
.W_7(W_7_x248),
.W_8(W_8_x248),
.W_9(W_9_x248)
) u_28X28_x248 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x248),
 .score_0 (score_0_x248),
 .score_1 (score_1_x248),
 .score_2 (score_2_x248),
 .score_3 (score_3_x248),
 .score_4 (score_4_x248),
 .score_5 (score_5_x248),
 .score_6 (score_6_x248),
 .score_7 (score_7_x248),
 .score_8 (score_8_x248),
 .score_9 (score_9_x248)
);
 
myram_28X28 #(
.ID(249),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x249),
.W_1(W_1_x249),
.W_2(W_2_x249),
.W_3(W_3_x249),
.W_4(W_4_x249),
.W_5(W_5_x249),
.W_6(W_6_x249),
.W_7(W_7_x249),
.W_8(W_8_x249),
.W_9(W_9_x249)
) u_28X28_x249 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x249),
 .score_0 (score_0_x249),
 .score_1 (score_1_x249),
 .score_2 (score_2_x249),
 .score_3 (score_3_x249),
 .score_4 (score_4_x249),
 .score_5 (score_5_x249),
 .score_6 (score_6_x249),
 .score_7 (score_7_x249),
 .score_8 (score_8_x249),
 .score_9 (score_9_x249)
);
 
myram_28X28 #(
.ID(250),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x250),
.W_1(W_1_x250),
.W_2(W_2_x250),
.W_3(W_3_x250),
.W_4(W_4_x250),
.W_5(W_5_x250),
.W_6(W_6_x250),
.W_7(W_7_x250),
.W_8(W_8_x250),
.W_9(W_9_x250)
) u_28X28_x250 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x250),
 .score_0 (score_0_x250),
 .score_1 (score_1_x250),
 .score_2 (score_2_x250),
 .score_3 (score_3_x250),
 .score_4 (score_4_x250),
 .score_5 (score_5_x250),
 .score_6 (score_6_x250),
 .score_7 (score_7_x250),
 .score_8 (score_8_x250),
 .score_9 (score_9_x250)
);
 
myram_28X28 #(
.ID(251),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x251),
.W_1(W_1_x251),
.W_2(W_2_x251),
.W_3(W_3_x251),
.W_4(W_4_x251),
.W_5(W_5_x251),
.W_6(W_6_x251),
.W_7(W_7_x251),
.W_8(W_8_x251),
.W_9(W_9_x251)
) u_28X28_x251 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x251),
 .score_0 (score_0_x251),
 .score_1 (score_1_x251),
 .score_2 (score_2_x251),
 .score_3 (score_3_x251),
 .score_4 (score_4_x251),
 .score_5 (score_5_x251),
 .score_6 (score_6_x251),
 .score_7 (score_7_x251),
 .score_8 (score_8_x251),
 .score_9 (score_9_x251)
);
 
myram_28X28 #(
.ID(252),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x252),
.W_1(W_1_x252),
.W_2(W_2_x252),
.W_3(W_3_x252),
.W_4(W_4_x252),
.W_5(W_5_x252),
.W_6(W_6_x252),
.W_7(W_7_x252),
.W_8(W_8_x252),
.W_9(W_9_x252)
) u_28X28_x252 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x252),
 .score_0 (score_0_x252),
 .score_1 (score_1_x252),
 .score_2 (score_2_x252),
 .score_3 (score_3_x252),
 .score_4 (score_4_x252),
 .score_5 (score_5_x252),
 .score_6 (score_6_x252),
 .score_7 (score_7_x252),
 .score_8 (score_8_x252),
 .score_9 (score_9_x252)
);
 
myram_28X28 #(
.ID(253),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x253),
.W_1(W_1_x253),
.W_2(W_2_x253),
.W_3(W_3_x253),
.W_4(W_4_x253),
.W_5(W_5_x253),
.W_6(W_6_x253),
.W_7(W_7_x253),
.W_8(W_8_x253),
.W_9(W_9_x253)
) u_28X28_x253 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x253),
 .score_0 (score_0_x253),
 .score_1 (score_1_x253),
 .score_2 (score_2_x253),
 .score_3 (score_3_x253),
 .score_4 (score_4_x253),
 .score_5 (score_5_x253),
 .score_6 (score_6_x253),
 .score_7 (score_7_x253),
 .score_8 (score_8_x253),
 .score_9 (score_9_x253)
);
 
myram_28X28 #(
.ID(254),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x254),
.W_1(W_1_x254),
.W_2(W_2_x254),
.W_3(W_3_x254),
.W_4(W_4_x254),
.W_5(W_5_x254),
.W_6(W_6_x254),
.W_7(W_7_x254),
.W_8(W_8_x254),
.W_9(W_9_x254)
) u_28X28_x254 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x254),
 .score_0 (score_0_x254),
 .score_1 (score_1_x254),
 .score_2 (score_2_x254),
 .score_3 (score_3_x254),
 .score_4 (score_4_x254),
 .score_5 (score_5_x254),
 .score_6 (score_6_x254),
 .score_7 (score_7_x254),
 .score_8 (score_8_x254),
 .score_9 (score_9_x254)
);
 
myram_28X28 #(
.ID(255),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x255),
.W_1(W_1_x255),
.W_2(W_2_x255),
.W_3(W_3_x255),
.W_4(W_4_x255),
.W_5(W_5_x255),
.W_6(W_6_x255),
.W_7(W_7_x255),
.W_8(W_8_x255),
.W_9(W_9_x255)
) u_28X28_x255 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x255),
 .score_0 (score_0_x255),
 .score_1 (score_1_x255),
 .score_2 (score_2_x255),
 .score_3 (score_3_x255),
 .score_4 (score_4_x255),
 .score_5 (score_5_x255),
 .score_6 (score_6_x255),
 .score_7 (score_7_x255),
 .score_8 (score_8_x255),
 .score_9 (score_9_x255)
);
 
myram_28X28 #(
.ID(256),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x256),
.W_1(W_1_x256),
.W_2(W_2_x256),
.W_3(W_3_x256),
.W_4(W_4_x256),
.W_5(W_5_x256),
.W_6(W_6_x256),
.W_7(W_7_x256),
.W_8(W_8_x256),
.W_9(W_9_x256)
) u_28X28_x256 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x256),
 .score_0 (score_0_x256),
 .score_1 (score_1_x256),
 .score_2 (score_2_x256),
 .score_3 (score_3_x256),
 .score_4 (score_4_x256),
 .score_5 (score_5_x256),
 .score_6 (score_6_x256),
 .score_7 (score_7_x256),
 .score_8 (score_8_x256),
 .score_9 (score_9_x256)
);
 
myram_28X28 #(
.ID(257),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x257),
.W_1(W_1_x257),
.W_2(W_2_x257),
.W_3(W_3_x257),
.W_4(W_4_x257),
.W_5(W_5_x257),
.W_6(W_6_x257),
.W_7(W_7_x257),
.W_8(W_8_x257),
.W_9(W_9_x257)
) u_28X28_x257 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x257),
 .score_0 (score_0_x257),
 .score_1 (score_1_x257),
 .score_2 (score_2_x257),
 .score_3 (score_3_x257),
 .score_4 (score_4_x257),
 .score_5 (score_5_x257),
 .score_6 (score_6_x257),
 .score_7 (score_7_x257),
 .score_8 (score_8_x257),
 .score_9 (score_9_x257)
);
 
myram_28X28 #(
.ID(258),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x258),
.W_1(W_1_x258),
.W_2(W_2_x258),
.W_3(W_3_x258),
.W_4(W_4_x258),
.W_5(W_5_x258),
.W_6(W_6_x258),
.W_7(W_7_x258),
.W_8(W_8_x258),
.W_9(W_9_x258)
) u_28X28_x258 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x258),
 .score_0 (score_0_x258),
 .score_1 (score_1_x258),
 .score_2 (score_2_x258),
 .score_3 (score_3_x258),
 .score_4 (score_4_x258),
 .score_5 (score_5_x258),
 .score_6 (score_6_x258),
 .score_7 (score_7_x258),
 .score_8 (score_8_x258),
 .score_9 (score_9_x258)
);
 
myram_28X28 #(
.ID(259),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x259),
.W_1(W_1_x259),
.W_2(W_2_x259),
.W_3(W_3_x259),
.W_4(W_4_x259),
.W_5(W_5_x259),
.W_6(W_6_x259),
.W_7(W_7_x259),
.W_8(W_8_x259),
.W_9(W_9_x259)
) u_28X28_x259 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x259),
 .score_0 (score_0_x259),
 .score_1 (score_1_x259),
 .score_2 (score_2_x259),
 .score_3 (score_3_x259),
 .score_4 (score_4_x259),
 .score_5 (score_5_x259),
 .score_6 (score_6_x259),
 .score_7 (score_7_x259),
 .score_8 (score_8_x259),
 .score_9 (score_9_x259)
);
 
myram_28X28 #(
.ID(260),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x260),
.W_1(W_1_x260),
.W_2(W_2_x260),
.W_3(W_3_x260),
.W_4(W_4_x260),
.W_5(W_5_x260),
.W_6(W_6_x260),
.W_7(W_7_x260),
.W_8(W_8_x260),
.W_9(W_9_x260)
) u_28X28_x260 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x260),
 .score_0 (score_0_x260),
 .score_1 (score_1_x260),
 .score_2 (score_2_x260),
 .score_3 (score_3_x260),
 .score_4 (score_4_x260),
 .score_5 (score_5_x260),
 .score_6 (score_6_x260),
 .score_7 (score_7_x260),
 .score_8 (score_8_x260),
 .score_9 (score_9_x260)
);
 
myram_28X28 #(
.ID(261),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x261),
.W_1(W_1_x261),
.W_2(W_2_x261),
.W_3(W_3_x261),
.W_4(W_4_x261),
.W_5(W_5_x261),
.W_6(W_6_x261),
.W_7(W_7_x261),
.W_8(W_8_x261),
.W_9(W_9_x261)
) u_28X28_x261 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x261),
 .score_0 (score_0_x261),
 .score_1 (score_1_x261),
 .score_2 (score_2_x261),
 .score_3 (score_3_x261),
 .score_4 (score_4_x261),
 .score_5 (score_5_x261),
 .score_6 (score_6_x261),
 .score_7 (score_7_x261),
 .score_8 (score_8_x261),
 .score_9 (score_9_x261)
);
 
myram_28X28 #(
.ID(262),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x262),
.W_1(W_1_x262),
.W_2(W_2_x262),
.W_3(W_3_x262),
.W_4(W_4_x262),
.W_5(W_5_x262),
.W_6(W_6_x262),
.W_7(W_7_x262),
.W_8(W_8_x262),
.W_9(W_9_x262)
) u_28X28_x262 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x262),
 .score_0 (score_0_x262),
 .score_1 (score_1_x262),
 .score_2 (score_2_x262),
 .score_3 (score_3_x262),
 .score_4 (score_4_x262),
 .score_5 (score_5_x262),
 .score_6 (score_6_x262),
 .score_7 (score_7_x262),
 .score_8 (score_8_x262),
 .score_9 (score_9_x262)
);
 
myram_28X28 #(
.ID(263),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x263),
.W_1(W_1_x263),
.W_2(W_2_x263),
.W_3(W_3_x263),
.W_4(W_4_x263),
.W_5(W_5_x263),
.W_6(W_6_x263),
.W_7(W_7_x263),
.W_8(W_8_x263),
.W_9(W_9_x263)
) u_28X28_x263 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x263),
 .score_0 (score_0_x263),
 .score_1 (score_1_x263),
 .score_2 (score_2_x263),
 .score_3 (score_3_x263),
 .score_4 (score_4_x263),
 .score_5 (score_5_x263),
 .score_6 (score_6_x263),
 .score_7 (score_7_x263),
 .score_8 (score_8_x263),
 .score_9 (score_9_x263)
);
 
myram_28X28 #(
.ID(264),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x264),
.W_1(W_1_x264),
.W_2(W_2_x264),
.W_3(W_3_x264),
.W_4(W_4_x264),
.W_5(W_5_x264),
.W_6(W_6_x264),
.W_7(W_7_x264),
.W_8(W_8_x264),
.W_9(W_9_x264)
) u_28X28_x264 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x264),
 .score_0 (score_0_x264),
 .score_1 (score_1_x264),
 .score_2 (score_2_x264),
 .score_3 (score_3_x264),
 .score_4 (score_4_x264),
 .score_5 (score_5_x264),
 .score_6 (score_6_x264),
 .score_7 (score_7_x264),
 .score_8 (score_8_x264),
 .score_9 (score_9_x264)
);
 
myram_28X28 #(
.ID(265),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x265),
.W_1(W_1_x265),
.W_2(W_2_x265),
.W_3(W_3_x265),
.W_4(W_4_x265),
.W_5(W_5_x265),
.W_6(W_6_x265),
.W_7(W_7_x265),
.W_8(W_8_x265),
.W_9(W_9_x265)
) u_28X28_x265 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x265),
 .score_0 (score_0_x265),
 .score_1 (score_1_x265),
 .score_2 (score_2_x265),
 .score_3 (score_3_x265),
 .score_4 (score_4_x265),
 .score_5 (score_5_x265),
 .score_6 (score_6_x265),
 .score_7 (score_7_x265),
 .score_8 (score_8_x265),
 .score_9 (score_9_x265)
);
 
myram_28X28 #(
.ID(266),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x266),
.W_1(W_1_x266),
.W_2(W_2_x266),
.W_3(W_3_x266),
.W_4(W_4_x266),
.W_5(W_5_x266),
.W_6(W_6_x266),
.W_7(W_7_x266),
.W_8(W_8_x266),
.W_9(W_9_x266)
) u_28X28_x266 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x266),
 .score_0 (score_0_x266),
 .score_1 (score_1_x266),
 .score_2 (score_2_x266),
 .score_3 (score_3_x266),
 .score_4 (score_4_x266),
 .score_5 (score_5_x266),
 .score_6 (score_6_x266),
 .score_7 (score_7_x266),
 .score_8 (score_8_x266),
 .score_9 (score_9_x266)
);
 
myram_28X28 #(
.ID(267),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x267),
.W_1(W_1_x267),
.W_2(W_2_x267),
.W_3(W_3_x267),
.W_4(W_4_x267),
.W_5(W_5_x267),
.W_6(W_6_x267),
.W_7(W_7_x267),
.W_8(W_8_x267),
.W_9(W_9_x267)
) u_28X28_x267 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x267),
 .score_0 (score_0_x267),
 .score_1 (score_1_x267),
 .score_2 (score_2_x267),
 .score_3 (score_3_x267),
 .score_4 (score_4_x267),
 .score_5 (score_5_x267),
 .score_6 (score_6_x267),
 .score_7 (score_7_x267),
 .score_8 (score_8_x267),
 .score_9 (score_9_x267)
);
 
myram_28X28 #(
.ID(268),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x268),
.W_1(W_1_x268),
.W_2(W_2_x268),
.W_3(W_3_x268),
.W_4(W_4_x268),
.W_5(W_5_x268),
.W_6(W_6_x268),
.W_7(W_7_x268),
.W_8(W_8_x268),
.W_9(W_9_x268)
) u_28X28_x268 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x268),
 .score_0 (score_0_x268),
 .score_1 (score_1_x268),
 .score_2 (score_2_x268),
 .score_3 (score_3_x268),
 .score_4 (score_4_x268),
 .score_5 (score_5_x268),
 .score_6 (score_6_x268),
 .score_7 (score_7_x268),
 .score_8 (score_8_x268),
 .score_9 (score_9_x268)
);
 
myram_28X28 #(
.ID(269),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x269),
.W_1(W_1_x269),
.W_2(W_2_x269),
.W_3(W_3_x269),
.W_4(W_4_x269),
.W_5(W_5_x269),
.W_6(W_6_x269),
.W_7(W_7_x269),
.W_8(W_8_x269),
.W_9(W_9_x269)
) u_28X28_x269 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x269),
 .score_0 (score_0_x269),
 .score_1 (score_1_x269),
 .score_2 (score_2_x269),
 .score_3 (score_3_x269),
 .score_4 (score_4_x269),
 .score_5 (score_5_x269),
 .score_6 (score_6_x269),
 .score_7 (score_7_x269),
 .score_8 (score_8_x269),
 .score_9 (score_9_x269)
);
 
myram_28X28 #(
.ID(270),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x270),
.W_1(W_1_x270),
.W_2(W_2_x270),
.W_3(W_3_x270),
.W_4(W_4_x270),
.W_5(W_5_x270),
.W_6(W_6_x270),
.W_7(W_7_x270),
.W_8(W_8_x270),
.W_9(W_9_x270)
) u_28X28_x270 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x270),
 .score_0 (score_0_x270),
 .score_1 (score_1_x270),
 .score_2 (score_2_x270),
 .score_3 (score_3_x270),
 .score_4 (score_4_x270),
 .score_5 (score_5_x270),
 .score_6 (score_6_x270),
 .score_7 (score_7_x270),
 .score_8 (score_8_x270),
 .score_9 (score_9_x270)
);
 
myram_28X28 #(
.ID(271),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x271),
.W_1(W_1_x271),
.W_2(W_2_x271),
.W_3(W_3_x271),
.W_4(W_4_x271),
.W_5(W_5_x271),
.W_6(W_6_x271),
.W_7(W_7_x271),
.W_8(W_8_x271),
.W_9(W_9_x271)
) u_28X28_x271 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x271),
 .score_0 (score_0_x271),
 .score_1 (score_1_x271),
 .score_2 (score_2_x271),
 .score_3 (score_3_x271),
 .score_4 (score_4_x271),
 .score_5 (score_5_x271),
 .score_6 (score_6_x271),
 .score_7 (score_7_x271),
 .score_8 (score_8_x271),
 .score_9 (score_9_x271)
);
 
myram_28X28 #(
.ID(272),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x272),
.W_1(W_1_x272),
.W_2(W_2_x272),
.W_3(W_3_x272),
.W_4(W_4_x272),
.W_5(W_5_x272),
.W_6(W_6_x272),
.W_7(W_7_x272),
.W_8(W_8_x272),
.W_9(W_9_x272)
) u_28X28_x272 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x272),
 .score_0 (score_0_x272),
 .score_1 (score_1_x272),
 .score_2 (score_2_x272),
 .score_3 (score_3_x272),
 .score_4 (score_4_x272),
 .score_5 (score_5_x272),
 .score_6 (score_6_x272),
 .score_7 (score_7_x272),
 .score_8 (score_8_x272),
 .score_9 (score_9_x272)
);
 
myram_28X28 #(
.ID(273),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x273),
.W_1(W_1_x273),
.W_2(W_2_x273),
.W_3(W_3_x273),
.W_4(W_4_x273),
.W_5(W_5_x273),
.W_6(W_6_x273),
.W_7(W_7_x273),
.W_8(W_8_x273),
.W_9(W_9_x273)
) u_28X28_x273 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x273),
 .score_0 (score_0_x273),
 .score_1 (score_1_x273),
 .score_2 (score_2_x273),
 .score_3 (score_3_x273),
 .score_4 (score_4_x273),
 .score_5 (score_5_x273),
 .score_6 (score_6_x273),
 .score_7 (score_7_x273),
 .score_8 (score_8_x273),
 .score_9 (score_9_x273)
);
 
myram_28X28 #(
.ID(274),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x274),
.W_1(W_1_x274),
.W_2(W_2_x274),
.W_3(W_3_x274),
.W_4(W_4_x274),
.W_5(W_5_x274),
.W_6(W_6_x274),
.W_7(W_7_x274),
.W_8(W_8_x274),
.W_9(W_9_x274)
) u_28X28_x274 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x274),
 .score_0 (score_0_x274),
 .score_1 (score_1_x274),
 .score_2 (score_2_x274),
 .score_3 (score_3_x274),
 .score_4 (score_4_x274),
 .score_5 (score_5_x274),
 .score_6 (score_6_x274),
 .score_7 (score_7_x274),
 .score_8 (score_8_x274),
 .score_9 (score_9_x274)
);
 
myram_28X28 #(
.ID(275),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x275),
.W_1(W_1_x275),
.W_2(W_2_x275),
.W_3(W_3_x275),
.W_4(W_4_x275),
.W_5(W_5_x275),
.W_6(W_6_x275),
.W_7(W_7_x275),
.W_8(W_8_x275),
.W_9(W_9_x275)
) u_28X28_x275 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x275),
 .score_0 (score_0_x275),
 .score_1 (score_1_x275),
 .score_2 (score_2_x275),
 .score_3 (score_3_x275),
 .score_4 (score_4_x275),
 .score_5 (score_5_x275),
 .score_6 (score_6_x275),
 .score_7 (score_7_x275),
 .score_8 (score_8_x275),
 .score_9 (score_9_x275)
);
 
myram_28X28 #(
.ID(276),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x276),
.W_1(W_1_x276),
.W_2(W_2_x276),
.W_3(W_3_x276),
.W_4(W_4_x276),
.W_5(W_5_x276),
.W_6(W_6_x276),
.W_7(W_7_x276),
.W_8(W_8_x276),
.W_9(W_9_x276)
) u_28X28_x276 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x276),
 .score_0 (score_0_x276),
 .score_1 (score_1_x276),
 .score_2 (score_2_x276),
 .score_3 (score_3_x276),
 .score_4 (score_4_x276),
 .score_5 (score_5_x276),
 .score_6 (score_6_x276),
 .score_7 (score_7_x276),
 .score_8 (score_8_x276),
 .score_9 (score_9_x276)
);
 
myram_28X28 #(
.ID(277),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x277),
.W_1(W_1_x277),
.W_2(W_2_x277),
.W_3(W_3_x277),
.W_4(W_4_x277),
.W_5(W_5_x277),
.W_6(W_6_x277),
.W_7(W_7_x277),
.W_8(W_8_x277),
.W_9(W_9_x277)
) u_28X28_x277 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x277),
 .score_0 (score_0_x277),
 .score_1 (score_1_x277),
 .score_2 (score_2_x277),
 .score_3 (score_3_x277),
 .score_4 (score_4_x277),
 .score_5 (score_5_x277),
 .score_6 (score_6_x277),
 .score_7 (score_7_x277),
 .score_8 (score_8_x277),
 .score_9 (score_9_x277)
);
 
myram_28X28 #(
.ID(278),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x278),
.W_1(W_1_x278),
.W_2(W_2_x278),
.W_3(W_3_x278),
.W_4(W_4_x278),
.W_5(W_5_x278),
.W_6(W_6_x278),
.W_7(W_7_x278),
.W_8(W_8_x278),
.W_9(W_9_x278)
) u_28X28_x278 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x278),
 .score_0 (score_0_x278),
 .score_1 (score_1_x278),
 .score_2 (score_2_x278),
 .score_3 (score_3_x278),
 .score_4 (score_4_x278),
 .score_5 (score_5_x278),
 .score_6 (score_6_x278),
 .score_7 (score_7_x278),
 .score_8 (score_8_x278),
 .score_9 (score_9_x278)
);
 
myram_28X28 #(
.ID(279),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x279),
.W_1(W_1_x279),
.W_2(W_2_x279),
.W_3(W_3_x279),
.W_4(W_4_x279),
.W_5(W_5_x279),
.W_6(W_6_x279),
.W_7(W_7_x279),
.W_8(W_8_x279),
.W_9(W_9_x279)
) u_28X28_x279 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x279),
 .score_0 (score_0_x279),
 .score_1 (score_1_x279),
 .score_2 (score_2_x279),
 .score_3 (score_3_x279),
 .score_4 (score_4_x279),
 .score_5 (score_5_x279),
 .score_6 (score_6_x279),
 .score_7 (score_7_x279),
 .score_8 (score_8_x279),
 .score_9 (score_9_x279)
);
 
myram_28X28 #(
.ID(280),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x280),
.W_1(W_1_x280),
.W_2(W_2_x280),
.W_3(W_3_x280),
.W_4(W_4_x280),
.W_5(W_5_x280),
.W_6(W_6_x280),
.W_7(W_7_x280),
.W_8(W_8_x280),
.W_9(W_9_x280)
) u_28X28_x280 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x280),
 .score_0 (score_0_x280),
 .score_1 (score_1_x280),
 .score_2 (score_2_x280),
 .score_3 (score_3_x280),
 .score_4 (score_4_x280),
 .score_5 (score_5_x280),
 .score_6 (score_6_x280),
 .score_7 (score_7_x280),
 .score_8 (score_8_x280),
 .score_9 (score_9_x280)
);
 
myram_28X28 #(
.ID(281),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x281),
.W_1(W_1_x281),
.W_2(W_2_x281),
.W_3(W_3_x281),
.W_4(W_4_x281),
.W_5(W_5_x281),
.W_6(W_6_x281),
.W_7(W_7_x281),
.W_8(W_8_x281),
.W_9(W_9_x281)
) u_28X28_x281 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x281),
 .score_0 (score_0_x281),
 .score_1 (score_1_x281),
 .score_2 (score_2_x281),
 .score_3 (score_3_x281),
 .score_4 (score_4_x281),
 .score_5 (score_5_x281),
 .score_6 (score_6_x281),
 .score_7 (score_7_x281),
 .score_8 (score_8_x281),
 .score_9 (score_9_x281)
);
 
myram_28X28 #(
.ID(282),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x282),
.W_1(W_1_x282),
.W_2(W_2_x282),
.W_3(W_3_x282),
.W_4(W_4_x282),
.W_5(W_5_x282),
.W_6(W_6_x282),
.W_7(W_7_x282),
.W_8(W_8_x282),
.W_9(W_9_x282)
) u_28X28_x282 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x282),
 .score_0 (score_0_x282),
 .score_1 (score_1_x282),
 .score_2 (score_2_x282),
 .score_3 (score_3_x282),
 .score_4 (score_4_x282),
 .score_5 (score_5_x282),
 .score_6 (score_6_x282),
 .score_7 (score_7_x282),
 .score_8 (score_8_x282),
 .score_9 (score_9_x282)
);
 
myram_28X28 #(
.ID(283),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x283),
.W_1(W_1_x283),
.W_2(W_2_x283),
.W_3(W_3_x283),
.W_4(W_4_x283),
.W_5(W_5_x283),
.W_6(W_6_x283),
.W_7(W_7_x283),
.W_8(W_8_x283),
.W_9(W_9_x283)
) u_28X28_x283 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x283),
 .score_0 (score_0_x283),
 .score_1 (score_1_x283),
 .score_2 (score_2_x283),
 .score_3 (score_3_x283),
 .score_4 (score_4_x283),
 .score_5 (score_5_x283),
 .score_6 (score_6_x283),
 .score_7 (score_7_x283),
 .score_8 (score_8_x283),
 .score_9 (score_9_x283)
);
 
myram_28X28 #(
.ID(284),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x284),
.W_1(W_1_x284),
.W_2(W_2_x284),
.W_3(W_3_x284),
.W_4(W_4_x284),
.W_5(W_5_x284),
.W_6(W_6_x284),
.W_7(W_7_x284),
.W_8(W_8_x284),
.W_9(W_9_x284)
) u_28X28_x284 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x284),
 .score_0 (score_0_x284),
 .score_1 (score_1_x284),
 .score_2 (score_2_x284),
 .score_3 (score_3_x284),
 .score_4 (score_4_x284),
 .score_5 (score_5_x284),
 .score_6 (score_6_x284),
 .score_7 (score_7_x284),
 .score_8 (score_8_x284),
 .score_9 (score_9_x284)
);
 
myram_28X28 #(
.ID(285),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x285),
.W_1(W_1_x285),
.W_2(W_2_x285),
.W_3(W_3_x285),
.W_4(W_4_x285),
.W_5(W_5_x285),
.W_6(W_6_x285),
.W_7(W_7_x285),
.W_8(W_8_x285),
.W_9(W_9_x285)
) u_28X28_x285 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x285),
 .score_0 (score_0_x285),
 .score_1 (score_1_x285),
 .score_2 (score_2_x285),
 .score_3 (score_3_x285),
 .score_4 (score_4_x285),
 .score_5 (score_5_x285),
 .score_6 (score_6_x285),
 .score_7 (score_7_x285),
 .score_8 (score_8_x285),
 .score_9 (score_9_x285)
);
 
myram_28X28 #(
.ID(286),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x286),
.W_1(W_1_x286),
.W_2(W_2_x286),
.W_3(W_3_x286),
.W_4(W_4_x286),
.W_5(W_5_x286),
.W_6(W_6_x286),
.W_7(W_7_x286),
.W_8(W_8_x286),
.W_9(W_9_x286)
) u_28X28_x286 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x286),
 .score_0 (score_0_x286),
 .score_1 (score_1_x286),
 .score_2 (score_2_x286),
 .score_3 (score_3_x286),
 .score_4 (score_4_x286),
 .score_5 (score_5_x286),
 .score_6 (score_6_x286),
 .score_7 (score_7_x286),
 .score_8 (score_8_x286),
 .score_9 (score_9_x286)
);
 
myram_28X28 #(
.ID(287),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x287),
.W_1(W_1_x287),
.W_2(W_2_x287),
.W_3(W_3_x287),
.W_4(W_4_x287),
.W_5(W_5_x287),
.W_6(W_6_x287),
.W_7(W_7_x287),
.W_8(W_8_x287),
.W_9(W_9_x287)
) u_28X28_x287 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x287),
 .score_0 (score_0_x287),
 .score_1 (score_1_x287),
 .score_2 (score_2_x287),
 .score_3 (score_3_x287),
 .score_4 (score_4_x287),
 .score_5 (score_5_x287),
 .score_6 (score_6_x287),
 .score_7 (score_7_x287),
 .score_8 (score_8_x287),
 .score_9 (score_9_x287)
);
 
myram_28X28 #(
.ID(288),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x288),
.W_1(W_1_x288),
.W_2(W_2_x288),
.W_3(W_3_x288),
.W_4(W_4_x288),
.W_5(W_5_x288),
.W_6(W_6_x288),
.W_7(W_7_x288),
.W_8(W_8_x288),
.W_9(W_9_x288)
) u_28X28_x288 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x288),
 .score_0 (score_0_x288),
 .score_1 (score_1_x288),
 .score_2 (score_2_x288),
 .score_3 (score_3_x288),
 .score_4 (score_4_x288),
 .score_5 (score_5_x288),
 .score_6 (score_6_x288),
 .score_7 (score_7_x288),
 .score_8 (score_8_x288),
 .score_9 (score_9_x288)
);
 
myram_28X28 #(
.ID(289),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x289),
.W_1(W_1_x289),
.W_2(W_2_x289),
.W_3(W_3_x289),
.W_4(W_4_x289),
.W_5(W_5_x289),
.W_6(W_6_x289),
.W_7(W_7_x289),
.W_8(W_8_x289),
.W_9(W_9_x289)
) u_28X28_x289 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x289),
 .score_0 (score_0_x289),
 .score_1 (score_1_x289),
 .score_2 (score_2_x289),
 .score_3 (score_3_x289),
 .score_4 (score_4_x289),
 .score_5 (score_5_x289),
 .score_6 (score_6_x289),
 .score_7 (score_7_x289),
 .score_8 (score_8_x289),
 .score_9 (score_9_x289)
);
 
myram_28X28 #(
.ID(290),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x290),
.W_1(W_1_x290),
.W_2(W_2_x290),
.W_3(W_3_x290),
.W_4(W_4_x290),
.W_5(W_5_x290),
.W_6(W_6_x290),
.W_7(W_7_x290),
.W_8(W_8_x290),
.W_9(W_9_x290)
) u_28X28_x290 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x290),
 .score_0 (score_0_x290),
 .score_1 (score_1_x290),
 .score_2 (score_2_x290),
 .score_3 (score_3_x290),
 .score_4 (score_4_x290),
 .score_5 (score_5_x290),
 .score_6 (score_6_x290),
 .score_7 (score_7_x290),
 .score_8 (score_8_x290),
 .score_9 (score_9_x290)
);
 
myram_28X28 #(
.ID(291),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x291),
.W_1(W_1_x291),
.W_2(W_2_x291),
.W_3(W_3_x291),
.W_4(W_4_x291),
.W_5(W_5_x291),
.W_6(W_6_x291),
.W_7(W_7_x291),
.W_8(W_8_x291),
.W_9(W_9_x291)
) u_28X28_x291 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x291),
 .score_0 (score_0_x291),
 .score_1 (score_1_x291),
 .score_2 (score_2_x291),
 .score_3 (score_3_x291),
 .score_4 (score_4_x291),
 .score_5 (score_5_x291),
 .score_6 (score_6_x291),
 .score_7 (score_7_x291),
 .score_8 (score_8_x291),
 .score_9 (score_9_x291)
);
 
myram_28X28 #(
.ID(292),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x292),
.W_1(W_1_x292),
.W_2(W_2_x292),
.W_3(W_3_x292),
.W_4(W_4_x292),
.W_5(W_5_x292),
.W_6(W_6_x292),
.W_7(W_7_x292),
.W_8(W_8_x292),
.W_9(W_9_x292)
) u_28X28_x292 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x292),
 .score_0 (score_0_x292),
 .score_1 (score_1_x292),
 .score_2 (score_2_x292),
 .score_3 (score_3_x292),
 .score_4 (score_4_x292),
 .score_5 (score_5_x292),
 .score_6 (score_6_x292),
 .score_7 (score_7_x292),
 .score_8 (score_8_x292),
 .score_9 (score_9_x292)
);
 
myram_28X28 #(
.ID(293),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x293),
.W_1(W_1_x293),
.W_2(W_2_x293),
.W_3(W_3_x293),
.W_4(W_4_x293),
.W_5(W_5_x293),
.W_6(W_6_x293),
.W_7(W_7_x293),
.W_8(W_8_x293),
.W_9(W_9_x293)
) u_28X28_x293 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x293),
 .score_0 (score_0_x293),
 .score_1 (score_1_x293),
 .score_2 (score_2_x293),
 .score_3 (score_3_x293),
 .score_4 (score_4_x293),
 .score_5 (score_5_x293),
 .score_6 (score_6_x293),
 .score_7 (score_7_x293),
 .score_8 (score_8_x293),
 .score_9 (score_9_x293)
);
 
myram_28X28 #(
.ID(294),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x294),
.W_1(W_1_x294),
.W_2(W_2_x294),
.W_3(W_3_x294),
.W_4(W_4_x294),
.W_5(W_5_x294),
.W_6(W_6_x294),
.W_7(W_7_x294),
.W_8(W_8_x294),
.W_9(W_9_x294)
) u_28X28_x294 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x294),
 .score_0 (score_0_x294),
 .score_1 (score_1_x294),
 .score_2 (score_2_x294),
 .score_3 (score_3_x294),
 .score_4 (score_4_x294),
 .score_5 (score_5_x294),
 .score_6 (score_6_x294),
 .score_7 (score_7_x294),
 .score_8 (score_8_x294),
 .score_9 (score_9_x294)
);
 
myram_28X28 #(
.ID(295),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x295),
.W_1(W_1_x295),
.W_2(W_2_x295),
.W_3(W_3_x295),
.W_4(W_4_x295),
.W_5(W_5_x295),
.W_6(W_6_x295),
.W_7(W_7_x295),
.W_8(W_8_x295),
.W_9(W_9_x295)
) u_28X28_x295 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x295),
 .score_0 (score_0_x295),
 .score_1 (score_1_x295),
 .score_2 (score_2_x295),
 .score_3 (score_3_x295),
 .score_4 (score_4_x295),
 .score_5 (score_5_x295),
 .score_6 (score_6_x295),
 .score_7 (score_7_x295),
 .score_8 (score_8_x295),
 .score_9 (score_9_x295)
);
 
myram_28X28 #(
.ID(296),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x296),
.W_1(W_1_x296),
.W_2(W_2_x296),
.W_3(W_3_x296),
.W_4(W_4_x296),
.W_5(W_5_x296),
.W_6(W_6_x296),
.W_7(W_7_x296),
.W_8(W_8_x296),
.W_9(W_9_x296)
) u_28X28_x296 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x296),
 .score_0 (score_0_x296),
 .score_1 (score_1_x296),
 .score_2 (score_2_x296),
 .score_3 (score_3_x296),
 .score_4 (score_4_x296),
 .score_5 (score_5_x296),
 .score_6 (score_6_x296),
 .score_7 (score_7_x296),
 .score_8 (score_8_x296),
 .score_9 (score_9_x296)
);
 
myram_28X28 #(
.ID(297),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x297),
.W_1(W_1_x297),
.W_2(W_2_x297),
.W_3(W_3_x297),
.W_4(W_4_x297),
.W_5(W_5_x297),
.W_6(W_6_x297),
.W_7(W_7_x297),
.W_8(W_8_x297),
.W_9(W_9_x297)
) u_28X28_x297 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x297),
 .score_0 (score_0_x297),
 .score_1 (score_1_x297),
 .score_2 (score_2_x297),
 .score_3 (score_3_x297),
 .score_4 (score_4_x297),
 .score_5 (score_5_x297),
 .score_6 (score_6_x297),
 .score_7 (score_7_x297),
 .score_8 (score_8_x297),
 .score_9 (score_9_x297)
);
 
myram_28X28 #(
.ID(298),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x298),
.W_1(W_1_x298),
.W_2(W_2_x298),
.W_3(W_3_x298),
.W_4(W_4_x298),
.W_5(W_5_x298),
.W_6(W_6_x298),
.W_7(W_7_x298),
.W_8(W_8_x298),
.W_9(W_9_x298)
) u_28X28_x298 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x298),
 .score_0 (score_0_x298),
 .score_1 (score_1_x298),
 .score_2 (score_2_x298),
 .score_3 (score_3_x298),
 .score_4 (score_4_x298),
 .score_5 (score_5_x298),
 .score_6 (score_6_x298),
 .score_7 (score_7_x298),
 .score_8 (score_8_x298),
 .score_9 (score_9_x298)
);
 
myram_28X28 #(
.ID(299),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x299),
.W_1(W_1_x299),
.W_2(W_2_x299),
.W_3(W_3_x299),
.W_4(W_4_x299),
.W_5(W_5_x299),
.W_6(W_6_x299),
.W_7(W_7_x299),
.W_8(W_8_x299),
.W_9(W_9_x299)
) u_28X28_x299 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x299),
 .score_0 (score_0_x299),
 .score_1 (score_1_x299),
 .score_2 (score_2_x299),
 .score_3 (score_3_x299),
 .score_4 (score_4_x299),
 .score_5 (score_5_x299),
 .score_6 (score_6_x299),
 .score_7 (score_7_x299),
 .score_8 (score_8_x299),
 .score_9 (score_9_x299)
);
 
myram_28X28 #(
.ID(300),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x300),
.W_1(W_1_x300),
.W_2(W_2_x300),
.W_3(W_3_x300),
.W_4(W_4_x300),
.W_5(W_5_x300),
.W_6(W_6_x300),
.W_7(W_7_x300),
.W_8(W_8_x300),
.W_9(W_9_x300)
) u_28X28_x300 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x300),
 .score_0 (score_0_x300),
 .score_1 (score_1_x300),
 .score_2 (score_2_x300),
 .score_3 (score_3_x300),
 .score_4 (score_4_x300),
 .score_5 (score_5_x300),
 .score_6 (score_6_x300),
 .score_7 (score_7_x300),
 .score_8 (score_8_x300),
 .score_9 (score_9_x300)
);
 
myram_28X28 #(
.ID(301),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x301),
.W_1(W_1_x301),
.W_2(W_2_x301),
.W_3(W_3_x301),
.W_4(W_4_x301),
.W_5(W_5_x301),
.W_6(W_6_x301),
.W_7(W_7_x301),
.W_8(W_8_x301),
.W_9(W_9_x301)
) u_28X28_x301 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x301),
 .score_0 (score_0_x301),
 .score_1 (score_1_x301),
 .score_2 (score_2_x301),
 .score_3 (score_3_x301),
 .score_4 (score_4_x301),
 .score_5 (score_5_x301),
 .score_6 (score_6_x301),
 .score_7 (score_7_x301),
 .score_8 (score_8_x301),
 .score_9 (score_9_x301)
);
 
myram_28X28 #(
.ID(302),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x302),
.W_1(W_1_x302),
.W_2(W_2_x302),
.W_3(W_3_x302),
.W_4(W_4_x302),
.W_5(W_5_x302),
.W_6(W_6_x302),
.W_7(W_7_x302),
.W_8(W_8_x302),
.W_9(W_9_x302)
) u_28X28_x302 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x302),
 .score_0 (score_0_x302),
 .score_1 (score_1_x302),
 .score_2 (score_2_x302),
 .score_3 (score_3_x302),
 .score_4 (score_4_x302),
 .score_5 (score_5_x302),
 .score_6 (score_6_x302),
 .score_7 (score_7_x302),
 .score_8 (score_8_x302),
 .score_9 (score_9_x302)
);
 
myram_28X28 #(
.ID(303),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x303),
.W_1(W_1_x303),
.W_2(W_2_x303),
.W_3(W_3_x303),
.W_4(W_4_x303),
.W_5(W_5_x303),
.W_6(W_6_x303),
.W_7(W_7_x303),
.W_8(W_8_x303),
.W_9(W_9_x303)
) u_28X28_x303 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x303),
 .score_0 (score_0_x303),
 .score_1 (score_1_x303),
 .score_2 (score_2_x303),
 .score_3 (score_3_x303),
 .score_4 (score_4_x303),
 .score_5 (score_5_x303),
 .score_6 (score_6_x303),
 .score_7 (score_7_x303),
 .score_8 (score_8_x303),
 .score_9 (score_9_x303)
);
 
myram_28X28 #(
.ID(304),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x304),
.W_1(W_1_x304),
.W_2(W_2_x304),
.W_3(W_3_x304),
.W_4(W_4_x304),
.W_5(W_5_x304),
.W_6(W_6_x304),
.W_7(W_7_x304),
.W_8(W_8_x304),
.W_9(W_9_x304)
) u_28X28_x304 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x304),
 .score_0 (score_0_x304),
 .score_1 (score_1_x304),
 .score_2 (score_2_x304),
 .score_3 (score_3_x304),
 .score_4 (score_4_x304),
 .score_5 (score_5_x304),
 .score_6 (score_6_x304),
 .score_7 (score_7_x304),
 .score_8 (score_8_x304),
 .score_9 (score_9_x304)
);
 
myram_28X28 #(
.ID(305),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x305),
.W_1(W_1_x305),
.W_2(W_2_x305),
.W_3(W_3_x305),
.W_4(W_4_x305),
.W_5(W_5_x305),
.W_6(W_6_x305),
.W_7(W_7_x305),
.W_8(W_8_x305),
.W_9(W_9_x305)
) u_28X28_x305 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x305),
 .score_0 (score_0_x305),
 .score_1 (score_1_x305),
 .score_2 (score_2_x305),
 .score_3 (score_3_x305),
 .score_4 (score_4_x305),
 .score_5 (score_5_x305),
 .score_6 (score_6_x305),
 .score_7 (score_7_x305),
 .score_8 (score_8_x305),
 .score_9 (score_9_x305)
);
 
myram_28X28 #(
.ID(306),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x306),
.W_1(W_1_x306),
.W_2(W_2_x306),
.W_3(W_3_x306),
.W_4(W_4_x306),
.W_5(W_5_x306),
.W_6(W_6_x306),
.W_7(W_7_x306),
.W_8(W_8_x306),
.W_9(W_9_x306)
) u_28X28_x306 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x306),
 .score_0 (score_0_x306),
 .score_1 (score_1_x306),
 .score_2 (score_2_x306),
 .score_3 (score_3_x306),
 .score_4 (score_4_x306),
 .score_5 (score_5_x306),
 .score_6 (score_6_x306),
 .score_7 (score_7_x306),
 .score_8 (score_8_x306),
 .score_9 (score_9_x306)
);
 
myram_28X28 #(
.ID(307),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x307),
.W_1(W_1_x307),
.W_2(W_2_x307),
.W_3(W_3_x307),
.W_4(W_4_x307),
.W_5(W_5_x307),
.W_6(W_6_x307),
.W_7(W_7_x307),
.W_8(W_8_x307),
.W_9(W_9_x307)
) u_28X28_x307 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x307),
 .score_0 (score_0_x307),
 .score_1 (score_1_x307),
 .score_2 (score_2_x307),
 .score_3 (score_3_x307),
 .score_4 (score_4_x307),
 .score_5 (score_5_x307),
 .score_6 (score_6_x307),
 .score_7 (score_7_x307),
 .score_8 (score_8_x307),
 .score_9 (score_9_x307)
);
 
myram_28X28 #(
.ID(308),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x308),
.W_1(W_1_x308),
.W_2(W_2_x308),
.W_3(W_3_x308),
.W_4(W_4_x308),
.W_5(W_5_x308),
.W_6(W_6_x308),
.W_7(W_7_x308),
.W_8(W_8_x308),
.W_9(W_9_x308)
) u_28X28_x308 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x308),
 .score_0 (score_0_x308),
 .score_1 (score_1_x308),
 .score_2 (score_2_x308),
 .score_3 (score_3_x308),
 .score_4 (score_4_x308),
 .score_5 (score_5_x308),
 .score_6 (score_6_x308),
 .score_7 (score_7_x308),
 .score_8 (score_8_x308),
 .score_9 (score_9_x308)
);
 
myram_28X28 #(
.ID(309),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x309),
.W_1(W_1_x309),
.W_2(W_2_x309),
.W_3(W_3_x309),
.W_4(W_4_x309),
.W_5(W_5_x309),
.W_6(W_6_x309),
.W_7(W_7_x309),
.W_8(W_8_x309),
.W_9(W_9_x309)
) u_28X28_x309 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x309),
 .score_0 (score_0_x309),
 .score_1 (score_1_x309),
 .score_2 (score_2_x309),
 .score_3 (score_3_x309),
 .score_4 (score_4_x309),
 .score_5 (score_5_x309),
 .score_6 (score_6_x309),
 .score_7 (score_7_x309),
 .score_8 (score_8_x309),
 .score_9 (score_9_x309)
);
 
myram_28X28 #(
.ID(310),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x310),
.W_1(W_1_x310),
.W_2(W_2_x310),
.W_3(W_3_x310),
.W_4(W_4_x310),
.W_5(W_5_x310),
.W_6(W_6_x310),
.W_7(W_7_x310),
.W_8(W_8_x310),
.W_9(W_9_x310)
) u_28X28_x310 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x310),
 .score_0 (score_0_x310),
 .score_1 (score_1_x310),
 .score_2 (score_2_x310),
 .score_3 (score_3_x310),
 .score_4 (score_4_x310),
 .score_5 (score_5_x310),
 .score_6 (score_6_x310),
 .score_7 (score_7_x310),
 .score_8 (score_8_x310),
 .score_9 (score_9_x310)
);
 
myram_28X28 #(
.ID(311),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x311),
.W_1(W_1_x311),
.W_2(W_2_x311),
.W_3(W_3_x311),
.W_4(W_4_x311),
.W_5(W_5_x311),
.W_6(W_6_x311),
.W_7(W_7_x311),
.W_8(W_8_x311),
.W_9(W_9_x311)
) u_28X28_x311 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x311),
 .score_0 (score_0_x311),
 .score_1 (score_1_x311),
 .score_2 (score_2_x311),
 .score_3 (score_3_x311),
 .score_4 (score_4_x311),
 .score_5 (score_5_x311),
 .score_6 (score_6_x311),
 .score_7 (score_7_x311),
 .score_8 (score_8_x311),
 .score_9 (score_9_x311)
);
 
myram_28X28 #(
.ID(312),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x312),
.W_1(W_1_x312),
.W_2(W_2_x312),
.W_3(W_3_x312),
.W_4(W_4_x312),
.W_5(W_5_x312),
.W_6(W_6_x312),
.W_7(W_7_x312),
.W_8(W_8_x312),
.W_9(W_9_x312)
) u_28X28_x312 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x312),
 .score_0 (score_0_x312),
 .score_1 (score_1_x312),
 .score_2 (score_2_x312),
 .score_3 (score_3_x312),
 .score_4 (score_4_x312),
 .score_5 (score_5_x312),
 .score_6 (score_6_x312),
 .score_7 (score_7_x312),
 .score_8 (score_8_x312),
 .score_9 (score_9_x312)
);
 
myram_28X28 #(
.ID(313),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x313),
.W_1(W_1_x313),
.W_2(W_2_x313),
.W_3(W_3_x313),
.W_4(W_4_x313),
.W_5(W_5_x313),
.W_6(W_6_x313),
.W_7(W_7_x313),
.W_8(W_8_x313),
.W_9(W_9_x313)
) u_28X28_x313 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x313),
 .score_0 (score_0_x313),
 .score_1 (score_1_x313),
 .score_2 (score_2_x313),
 .score_3 (score_3_x313),
 .score_4 (score_4_x313),
 .score_5 (score_5_x313),
 .score_6 (score_6_x313),
 .score_7 (score_7_x313),
 .score_8 (score_8_x313),
 .score_9 (score_9_x313)
);
 
myram_28X28 #(
.ID(314),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x314),
.W_1(W_1_x314),
.W_2(W_2_x314),
.W_3(W_3_x314),
.W_4(W_4_x314),
.W_5(W_5_x314),
.W_6(W_6_x314),
.W_7(W_7_x314),
.W_8(W_8_x314),
.W_9(W_9_x314)
) u_28X28_x314 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x314),
 .score_0 (score_0_x314),
 .score_1 (score_1_x314),
 .score_2 (score_2_x314),
 .score_3 (score_3_x314),
 .score_4 (score_4_x314),
 .score_5 (score_5_x314),
 .score_6 (score_6_x314),
 .score_7 (score_7_x314),
 .score_8 (score_8_x314),
 .score_9 (score_9_x314)
);
 
myram_28X28 #(
.ID(315),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x315),
.W_1(W_1_x315),
.W_2(W_2_x315),
.W_3(W_3_x315),
.W_4(W_4_x315),
.W_5(W_5_x315),
.W_6(W_6_x315),
.W_7(W_7_x315),
.W_8(W_8_x315),
.W_9(W_9_x315)
) u_28X28_x315 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x315),
 .score_0 (score_0_x315),
 .score_1 (score_1_x315),
 .score_2 (score_2_x315),
 .score_3 (score_3_x315),
 .score_4 (score_4_x315),
 .score_5 (score_5_x315),
 .score_6 (score_6_x315),
 .score_7 (score_7_x315),
 .score_8 (score_8_x315),
 .score_9 (score_9_x315)
);
 
myram_28X28 #(
.ID(316),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x316),
.W_1(W_1_x316),
.W_2(W_2_x316),
.W_3(W_3_x316),
.W_4(W_4_x316),
.W_5(W_5_x316),
.W_6(W_6_x316),
.W_7(W_7_x316),
.W_8(W_8_x316),
.W_9(W_9_x316)
) u_28X28_x316 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x316),
 .score_0 (score_0_x316),
 .score_1 (score_1_x316),
 .score_2 (score_2_x316),
 .score_3 (score_3_x316),
 .score_4 (score_4_x316),
 .score_5 (score_5_x316),
 .score_6 (score_6_x316),
 .score_7 (score_7_x316),
 .score_8 (score_8_x316),
 .score_9 (score_9_x316)
);
 
myram_28X28 #(
.ID(317),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x317),
.W_1(W_1_x317),
.W_2(W_2_x317),
.W_3(W_3_x317),
.W_4(W_4_x317),
.W_5(W_5_x317),
.W_6(W_6_x317),
.W_7(W_7_x317),
.W_8(W_8_x317),
.W_9(W_9_x317)
) u_28X28_x317 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x317),
 .score_0 (score_0_x317),
 .score_1 (score_1_x317),
 .score_2 (score_2_x317),
 .score_3 (score_3_x317),
 .score_4 (score_4_x317),
 .score_5 (score_5_x317),
 .score_6 (score_6_x317),
 .score_7 (score_7_x317),
 .score_8 (score_8_x317),
 .score_9 (score_9_x317)
);
 
myram_28X28 #(
.ID(318),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x318),
.W_1(W_1_x318),
.W_2(W_2_x318),
.W_3(W_3_x318),
.W_4(W_4_x318),
.W_5(W_5_x318),
.W_6(W_6_x318),
.W_7(W_7_x318),
.W_8(W_8_x318),
.W_9(W_9_x318)
) u_28X28_x318 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x318),
 .score_0 (score_0_x318),
 .score_1 (score_1_x318),
 .score_2 (score_2_x318),
 .score_3 (score_3_x318),
 .score_4 (score_4_x318),
 .score_5 (score_5_x318),
 .score_6 (score_6_x318),
 .score_7 (score_7_x318),
 .score_8 (score_8_x318),
 .score_9 (score_9_x318)
);
 
myram_28X28 #(
.ID(319),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x319),
.W_1(W_1_x319),
.W_2(W_2_x319),
.W_3(W_3_x319),
.W_4(W_4_x319),
.W_5(W_5_x319),
.W_6(W_6_x319),
.W_7(W_7_x319),
.W_8(W_8_x319),
.W_9(W_9_x319)
) u_28X28_x319 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x319),
 .score_0 (score_0_x319),
 .score_1 (score_1_x319),
 .score_2 (score_2_x319),
 .score_3 (score_3_x319),
 .score_4 (score_4_x319),
 .score_5 (score_5_x319),
 .score_6 (score_6_x319),
 .score_7 (score_7_x319),
 .score_8 (score_8_x319),
 .score_9 (score_9_x319)
);
 
myram_28X28 #(
.ID(320),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x320),
.W_1(W_1_x320),
.W_2(W_2_x320),
.W_3(W_3_x320),
.W_4(W_4_x320),
.W_5(W_5_x320),
.W_6(W_6_x320),
.W_7(W_7_x320),
.W_8(W_8_x320),
.W_9(W_9_x320)
) u_28X28_x320 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x320),
 .score_0 (score_0_x320),
 .score_1 (score_1_x320),
 .score_2 (score_2_x320),
 .score_3 (score_3_x320),
 .score_4 (score_4_x320),
 .score_5 (score_5_x320),
 .score_6 (score_6_x320),
 .score_7 (score_7_x320),
 .score_8 (score_8_x320),
 .score_9 (score_9_x320)
);
 
myram_28X28 #(
.ID(321),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x321),
.W_1(W_1_x321),
.W_2(W_2_x321),
.W_3(W_3_x321),
.W_4(W_4_x321),
.W_5(W_5_x321),
.W_6(W_6_x321),
.W_7(W_7_x321),
.W_8(W_8_x321),
.W_9(W_9_x321)
) u_28X28_x321 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x321),
 .score_0 (score_0_x321),
 .score_1 (score_1_x321),
 .score_2 (score_2_x321),
 .score_3 (score_3_x321),
 .score_4 (score_4_x321),
 .score_5 (score_5_x321),
 .score_6 (score_6_x321),
 .score_7 (score_7_x321),
 .score_8 (score_8_x321),
 .score_9 (score_9_x321)
);
 
myram_28X28 #(
.ID(322),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x322),
.W_1(W_1_x322),
.W_2(W_2_x322),
.W_3(W_3_x322),
.W_4(W_4_x322),
.W_5(W_5_x322),
.W_6(W_6_x322),
.W_7(W_7_x322),
.W_8(W_8_x322),
.W_9(W_9_x322)
) u_28X28_x322 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x322),
 .score_0 (score_0_x322),
 .score_1 (score_1_x322),
 .score_2 (score_2_x322),
 .score_3 (score_3_x322),
 .score_4 (score_4_x322),
 .score_5 (score_5_x322),
 .score_6 (score_6_x322),
 .score_7 (score_7_x322),
 .score_8 (score_8_x322),
 .score_9 (score_9_x322)
);
 
myram_28X28 #(
.ID(323),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x323),
.W_1(W_1_x323),
.W_2(W_2_x323),
.W_3(W_3_x323),
.W_4(W_4_x323),
.W_5(W_5_x323),
.W_6(W_6_x323),
.W_7(W_7_x323),
.W_8(W_8_x323),
.W_9(W_9_x323)
) u_28X28_x323 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x323),
 .score_0 (score_0_x323),
 .score_1 (score_1_x323),
 .score_2 (score_2_x323),
 .score_3 (score_3_x323),
 .score_4 (score_4_x323),
 .score_5 (score_5_x323),
 .score_6 (score_6_x323),
 .score_7 (score_7_x323),
 .score_8 (score_8_x323),
 .score_9 (score_9_x323)
);
 
myram_28X28 #(
.ID(324),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x324),
.W_1(W_1_x324),
.W_2(W_2_x324),
.W_3(W_3_x324),
.W_4(W_4_x324),
.W_5(W_5_x324),
.W_6(W_6_x324),
.W_7(W_7_x324),
.W_8(W_8_x324),
.W_9(W_9_x324)
) u_28X28_x324 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x324),
 .score_0 (score_0_x324),
 .score_1 (score_1_x324),
 .score_2 (score_2_x324),
 .score_3 (score_3_x324),
 .score_4 (score_4_x324),
 .score_5 (score_5_x324),
 .score_6 (score_6_x324),
 .score_7 (score_7_x324),
 .score_8 (score_8_x324),
 .score_9 (score_9_x324)
);
 
myram_28X28 #(
.ID(325),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x325),
.W_1(W_1_x325),
.W_2(W_2_x325),
.W_3(W_3_x325),
.W_4(W_4_x325),
.W_5(W_5_x325),
.W_6(W_6_x325),
.W_7(W_7_x325),
.W_8(W_8_x325),
.W_9(W_9_x325)
) u_28X28_x325 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x325),
 .score_0 (score_0_x325),
 .score_1 (score_1_x325),
 .score_2 (score_2_x325),
 .score_3 (score_3_x325),
 .score_4 (score_4_x325),
 .score_5 (score_5_x325),
 .score_6 (score_6_x325),
 .score_7 (score_7_x325),
 .score_8 (score_8_x325),
 .score_9 (score_9_x325)
);
 
myram_28X28 #(
.ID(326),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x326),
.W_1(W_1_x326),
.W_2(W_2_x326),
.W_3(W_3_x326),
.W_4(W_4_x326),
.W_5(W_5_x326),
.W_6(W_6_x326),
.W_7(W_7_x326),
.W_8(W_8_x326),
.W_9(W_9_x326)
) u_28X28_x326 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x326),
 .score_0 (score_0_x326),
 .score_1 (score_1_x326),
 .score_2 (score_2_x326),
 .score_3 (score_3_x326),
 .score_4 (score_4_x326),
 .score_5 (score_5_x326),
 .score_6 (score_6_x326),
 .score_7 (score_7_x326),
 .score_8 (score_8_x326),
 .score_9 (score_9_x326)
);
 
myram_28X28 #(
.ID(327),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x327),
.W_1(W_1_x327),
.W_2(W_2_x327),
.W_3(W_3_x327),
.W_4(W_4_x327),
.W_5(W_5_x327),
.W_6(W_6_x327),
.W_7(W_7_x327),
.W_8(W_8_x327),
.W_9(W_9_x327)
) u_28X28_x327 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x327),
 .score_0 (score_0_x327),
 .score_1 (score_1_x327),
 .score_2 (score_2_x327),
 .score_3 (score_3_x327),
 .score_4 (score_4_x327),
 .score_5 (score_5_x327),
 .score_6 (score_6_x327),
 .score_7 (score_7_x327),
 .score_8 (score_8_x327),
 .score_9 (score_9_x327)
);
 
myram_28X28 #(
.ID(328),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x328),
.W_1(W_1_x328),
.W_2(W_2_x328),
.W_3(W_3_x328),
.W_4(W_4_x328),
.W_5(W_5_x328),
.W_6(W_6_x328),
.W_7(W_7_x328),
.W_8(W_8_x328),
.W_9(W_9_x328)
) u_28X28_x328 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x328),
 .score_0 (score_0_x328),
 .score_1 (score_1_x328),
 .score_2 (score_2_x328),
 .score_3 (score_3_x328),
 .score_4 (score_4_x328),
 .score_5 (score_5_x328),
 .score_6 (score_6_x328),
 .score_7 (score_7_x328),
 .score_8 (score_8_x328),
 .score_9 (score_9_x328)
);
 
myram_28X28 #(
.ID(329),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x329),
.W_1(W_1_x329),
.W_2(W_2_x329),
.W_3(W_3_x329),
.W_4(W_4_x329),
.W_5(W_5_x329),
.W_6(W_6_x329),
.W_7(W_7_x329),
.W_8(W_8_x329),
.W_9(W_9_x329)
) u_28X28_x329 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x329),
 .score_0 (score_0_x329),
 .score_1 (score_1_x329),
 .score_2 (score_2_x329),
 .score_3 (score_3_x329),
 .score_4 (score_4_x329),
 .score_5 (score_5_x329),
 .score_6 (score_6_x329),
 .score_7 (score_7_x329),
 .score_8 (score_8_x329),
 .score_9 (score_9_x329)
);
 
myram_28X28 #(
.ID(330),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x330),
.W_1(W_1_x330),
.W_2(W_2_x330),
.W_3(W_3_x330),
.W_4(W_4_x330),
.W_5(W_5_x330),
.W_6(W_6_x330),
.W_7(W_7_x330),
.W_8(W_8_x330),
.W_9(W_9_x330)
) u_28X28_x330 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x330),
 .score_0 (score_0_x330),
 .score_1 (score_1_x330),
 .score_2 (score_2_x330),
 .score_3 (score_3_x330),
 .score_4 (score_4_x330),
 .score_5 (score_5_x330),
 .score_6 (score_6_x330),
 .score_7 (score_7_x330),
 .score_8 (score_8_x330),
 .score_9 (score_9_x330)
);
 
myram_28X28 #(
.ID(331),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x331),
.W_1(W_1_x331),
.W_2(W_2_x331),
.W_3(W_3_x331),
.W_4(W_4_x331),
.W_5(W_5_x331),
.W_6(W_6_x331),
.W_7(W_7_x331),
.W_8(W_8_x331),
.W_9(W_9_x331)
) u_28X28_x331 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x331),
 .score_0 (score_0_x331),
 .score_1 (score_1_x331),
 .score_2 (score_2_x331),
 .score_3 (score_3_x331),
 .score_4 (score_4_x331),
 .score_5 (score_5_x331),
 .score_6 (score_6_x331),
 .score_7 (score_7_x331),
 .score_8 (score_8_x331),
 .score_9 (score_9_x331)
);
 
myram_28X28 #(
.ID(332),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x332),
.W_1(W_1_x332),
.W_2(W_2_x332),
.W_3(W_3_x332),
.W_4(W_4_x332),
.W_5(W_5_x332),
.W_6(W_6_x332),
.W_7(W_7_x332),
.W_8(W_8_x332),
.W_9(W_9_x332)
) u_28X28_x332 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x332),
 .score_0 (score_0_x332),
 .score_1 (score_1_x332),
 .score_2 (score_2_x332),
 .score_3 (score_3_x332),
 .score_4 (score_4_x332),
 .score_5 (score_5_x332),
 .score_6 (score_6_x332),
 .score_7 (score_7_x332),
 .score_8 (score_8_x332),
 .score_9 (score_9_x332)
);
 
myram_28X28 #(
.ID(333),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x333),
.W_1(W_1_x333),
.W_2(W_2_x333),
.W_3(W_3_x333),
.W_4(W_4_x333),
.W_5(W_5_x333),
.W_6(W_6_x333),
.W_7(W_7_x333),
.W_8(W_8_x333),
.W_9(W_9_x333)
) u_28X28_x333 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x333),
 .score_0 (score_0_x333),
 .score_1 (score_1_x333),
 .score_2 (score_2_x333),
 .score_3 (score_3_x333),
 .score_4 (score_4_x333),
 .score_5 (score_5_x333),
 .score_6 (score_6_x333),
 .score_7 (score_7_x333),
 .score_8 (score_8_x333),
 .score_9 (score_9_x333)
);
 
myram_28X28 #(
.ID(334),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x334),
.W_1(W_1_x334),
.W_2(W_2_x334),
.W_3(W_3_x334),
.W_4(W_4_x334),
.W_5(W_5_x334),
.W_6(W_6_x334),
.W_7(W_7_x334),
.W_8(W_8_x334),
.W_9(W_9_x334)
) u_28X28_x334 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x334),
 .score_0 (score_0_x334),
 .score_1 (score_1_x334),
 .score_2 (score_2_x334),
 .score_3 (score_3_x334),
 .score_4 (score_4_x334),
 .score_5 (score_5_x334),
 .score_6 (score_6_x334),
 .score_7 (score_7_x334),
 .score_8 (score_8_x334),
 .score_9 (score_9_x334)
);
 
myram_28X28 #(
.ID(335),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x335),
.W_1(W_1_x335),
.W_2(W_2_x335),
.W_3(W_3_x335),
.W_4(W_4_x335),
.W_5(W_5_x335),
.W_6(W_6_x335),
.W_7(W_7_x335),
.W_8(W_8_x335),
.W_9(W_9_x335)
) u_28X28_x335 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x335),
 .score_0 (score_0_x335),
 .score_1 (score_1_x335),
 .score_2 (score_2_x335),
 .score_3 (score_3_x335),
 .score_4 (score_4_x335),
 .score_5 (score_5_x335),
 .score_6 (score_6_x335),
 .score_7 (score_7_x335),
 .score_8 (score_8_x335),
 .score_9 (score_9_x335)
);
 
myram_28X28 #(
.ID(336),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x336),
.W_1(W_1_x336),
.W_2(W_2_x336),
.W_3(W_3_x336),
.W_4(W_4_x336),
.W_5(W_5_x336),
.W_6(W_6_x336),
.W_7(W_7_x336),
.W_8(W_8_x336),
.W_9(W_9_x336)
) u_28X28_x336 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x336),
 .score_0 (score_0_x336),
 .score_1 (score_1_x336),
 .score_2 (score_2_x336),
 .score_3 (score_3_x336),
 .score_4 (score_4_x336),
 .score_5 (score_5_x336),
 .score_6 (score_6_x336),
 .score_7 (score_7_x336),
 .score_8 (score_8_x336),
 .score_9 (score_9_x336)
);
 
myram_28X28 #(
.ID(337),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x337),
.W_1(W_1_x337),
.W_2(W_2_x337),
.W_3(W_3_x337),
.W_4(W_4_x337),
.W_5(W_5_x337),
.W_6(W_6_x337),
.W_7(W_7_x337),
.W_8(W_8_x337),
.W_9(W_9_x337)
) u_28X28_x337 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x337),
 .score_0 (score_0_x337),
 .score_1 (score_1_x337),
 .score_2 (score_2_x337),
 .score_3 (score_3_x337),
 .score_4 (score_4_x337),
 .score_5 (score_5_x337),
 .score_6 (score_6_x337),
 .score_7 (score_7_x337),
 .score_8 (score_8_x337),
 .score_9 (score_9_x337)
);
 
myram_28X28 #(
.ID(338),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x338),
.W_1(W_1_x338),
.W_2(W_2_x338),
.W_3(W_3_x338),
.W_4(W_4_x338),
.W_5(W_5_x338),
.W_6(W_6_x338),
.W_7(W_7_x338),
.W_8(W_8_x338),
.W_9(W_9_x338)
) u_28X28_x338 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x338),
 .score_0 (score_0_x338),
 .score_1 (score_1_x338),
 .score_2 (score_2_x338),
 .score_3 (score_3_x338),
 .score_4 (score_4_x338),
 .score_5 (score_5_x338),
 .score_6 (score_6_x338),
 .score_7 (score_7_x338),
 .score_8 (score_8_x338),
 .score_9 (score_9_x338)
);
 
myram_28X28 #(
.ID(339),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x339),
.W_1(W_1_x339),
.W_2(W_2_x339),
.W_3(W_3_x339),
.W_4(W_4_x339),
.W_5(W_5_x339),
.W_6(W_6_x339),
.W_7(W_7_x339),
.W_8(W_8_x339),
.W_9(W_9_x339)
) u_28X28_x339 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x339),
 .score_0 (score_0_x339),
 .score_1 (score_1_x339),
 .score_2 (score_2_x339),
 .score_3 (score_3_x339),
 .score_4 (score_4_x339),
 .score_5 (score_5_x339),
 .score_6 (score_6_x339),
 .score_7 (score_7_x339),
 .score_8 (score_8_x339),
 .score_9 (score_9_x339)
);
 
myram_28X28 #(
.ID(340),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x340),
.W_1(W_1_x340),
.W_2(W_2_x340),
.W_3(W_3_x340),
.W_4(W_4_x340),
.W_5(W_5_x340),
.W_6(W_6_x340),
.W_7(W_7_x340),
.W_8(W_8_x340),
.W_9(W_9_x340)
) u_28X28_x340 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x340),
 .score_0 (score_0_x340),
 .score_1 (score_1_x340),
 .score_2 (score_2_x340),
 .score_3 (score_3_x340),
 .score_4 (score_4_x340),
 .score_5 (score_5_x340),
 .score_6 (score_6_x340),
 .score_7 (score_7_x340),
 .score_8 (score_8_x340),
 .score_9 (score_9_x340)
);
 
myram_28X28 #(
.ID(341),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x341),
.W_1(W_1_x341),
.W_2(W_2_x341),
.W_3(W_3_x341),
.W_4(W_4_x341),
.W_5(W_5_x341),
.W_6(W_6_x341),
.W_7(W_7_x341),
.W_8(W_8_x341),
.W_9(W_9_x341)
) u_28X28_x341 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x341),
 .score_0 (score_0_x341),
 .score_1 (score_1_x341),
 .score_2 (score_2_x341),
 .score_3 (score_3_x341),
 .score_4 (score_4_x341),
 .score_5 (score_5_x341),
 .score_6 (score_6_x341),
 .score_7 (score_7_x341),
 .score_8 (score_8_x341),
 .score_9 (score_9_x341)
);
 
myram_28X28 #(
.ID(342),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x342),
.W_1(W_1_x342),
.W_2(W_2_x342),
.W_3(W_3_x342),
.W_4(W_4_x342),
.W_5(W_5_x342),
.W_6(W_6_x342),
.W_7(W_7_x342),
.W_8(W_8_x342),
.W_9(W_9_x342)
) u_28X28_x342 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x342),
 .score_0 (score_0_x342),
 .score_1 (score_1_x342),
 .score_2 (score_2_x342),
 .score_3 (score_3_x342),
 .score_4 (score_4_x342),
 .score_5 (score_5_x342),
 .score_6 (score_6_x342),
 .score_7 (score_7_x342),
 .score_8 (score_8_x342),
 .score_9 (score_9_x342)
);
 
myram_28X28 #(
.ID(343),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x343),
.W_1(W_1_x343),
.W_2(W_2_x343),
.W_3(W_3_x343),
.W_4(W_4_x343),
.W_5(W_5_x343),
.W_6(W_6_x343),
.W_7(W_7_x343),
.W_8(W_8_x343),
.W_9(W_9_x343)
) u_28X28_x343 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x343),
 .score_0 (score_0_x343),
 .score_1 (score_1_x343),
 .score_2 (score_2_x343),
 .score_3 (score_3_x343),
 .score_4 (score_4_x343),
 .score_5 (score_5_x343),
 .score_6 (score_6_x343),
 .score_7 (score_7_x343),
 .score_8 (score_8_x343),
 .score_9 (score_9_x343)
);
 
myram_28X28 #(
.ID(344),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x344),
.W_1(W_1_x344),
.W_2(W_2_x344),
.W_3(W_3_x344),
.W_4(W_4_x344),
.W_5(W_5_x344),
.W_6(W_6_x344),
.W_7(W_7_x344),
.W_8(W_8_x344),
.W_9(W_9_x344)
) u_28X28_x344 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x344),
 .score_0 (score_0_x344),
 .score_1 (score_1_x344),
 .score_2 (score_2_x344),
 .score_3 (score_3_x344),
 .score_4 (score_4_x344),
 .score_5 (score_5_x344),
 .score_6 (score_6_x344),
 .score_7 (score_7_x344),
 .score_8 (score_8_x344),
 .score_9 (score_9_x344)
);
 
myram_28X28 #(
.ID(345),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x345),
.W_1(W_1_x345),
.W_2(W_2_x345),
.W_3(W_3_x345),
.W_4(W_4_x345),
.W_5(W_5_x345),
.W_6(W_6_x345),
.W_7(W_7_x345),
.W_8(W_8_x345),
.W_9(W_9_x345)
) u_28X28_x345 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x345),
 .score_0 (score_0_x345),
 .score_1 (score_1_x345),
 .score_2 (score_2_x345),
 .score_3 (score_3_x345),
 .score_4 (score_4_x345),
 .score_5 (score_5_x345),
 .score_6 (score_6_x345),
 .score_7 (score_7_x345),
 .score_8 (score_8_x345),
 .score_9 (score_9_x345)
);
 
myram_28X28 #(
.ID(346),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x346),
.W_1(W_1_x346),
.W_2(W_2_x346),
.W_3(W_3_x346),
.W_4(W_4_x346),
.W_5(W_5_x346),
.W_6(W_6_x346),
.W_7(W_7_x346),
.W_8(W_8_x346),
.W_9(W_9_x346)
) u_28X28_x346 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x346),
 .score_0 (score_0_x346),
 .score_1 (score_1_x346),
 .score_2 (score_2_x346),
 .score_3 (score_3_x346),
 .score_4 (score_4_x346),
 .score_5 (score_5_x346),
 .score_6 (score_6_x346),
 .score_7 (score_7_x346),
 .score_8 (score_8_x346),
 .score_9 (score_9_x346)
);
 
myram_28X28 #(
.ID(347),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x347),
.W_1(W_1_x347),
.W_2(W_2_x347),
.W_3(W_3_x347),
.W_4(W_4_x347),
.W_5(W_5_x347),
.W_6(W_6_x347),
.W_7(W_7_x347),
.W_8(W_8_x347),
.W_9(W_9_x347)
) u_28X28_x347 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x347),
 .score_0 (score_0_x347),
 .score_1 (score_1_x347),
 .score_2 (score_2_x347),
 .score_3 (score_3_x347),
 .score_4 (score_4_x347),
 .score_5 (score_5_x347),
 .score_6 (score_6_x347),
 .score_7 (score_7_x347),
 .score_8 (score_8_x347),
 .score_9 (score_9_x347)
);
 
myram_28X28 #(
.ID(348),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x348),
.W_1(W_1_x348),
.W_2(W_2_x348),
.W_3(W_3_x348),
.W_4(W_4_x348),
.W_5(W_5_x348),
.W_6(W_6_x348),
.W_7(W_7_x348),
.W_8(W_8_x348),
.W_9(W_9_x348)
) u_28X28_x348 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x348),
 .score_0 (score_0_x348),
 .score_1 (score_1_x348),
 .score_2 (score_2_x348),
 .score_3 (score_3_x348),
 .score_4 (score_4_x348),
 .score_5 (score_5_x348),
 .score_6 (score_6_x348),
 .score_7 (score_7_x348),
 .score_8 (score_8_x348),
 .score_9 (score_9_x348)
);
 
myram_28X28 #(
.ID(349),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x349),
.W_1(W_1_x349),
.W_2(W_2_x349),
.W_3(W_3_x349),
.W_4(W_4_x349),
.W_5(W_5_x349),
.W_6(W_6_x349),
.W_7(W_7_x349),
.W_8(W_8_x349),
.W_9(W_9_x349)
) u_28X28_x349 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x349),
 .score_0 (score_0_x349),
 .score_1 (score_1_x349),
 .score_2 (score_2_x349),
 .score_3 (score_3_x349),
 .score_4 (score_4_x349),
 .score_5 (score_5_x349),
 .score_6 (score_6_x349),
 .score_7 (score_7_x349),
 .score_8 (score_8_x349),
 .score_9 (score_9_x349)
);
 
myram_28X28 #(
.ID(350),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x350),
.W_1(W_1_x350),
.W_2(W_2_x350),
.W_3(W_3_x350),
.W_4(W_4_x350),
.W_5(W_5_x350),
.W_6(W_6_x350),
.W_7(W_7_x350),
.W_8(W_8_x350),
.W_9(W_9_x350)
) u_28X28_x350 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x350),
 .score_0 (score_0_x350),
 .score_1 (score_1_x350),
 .score_2 (score_2_x350),
 .score_3 (score_3_x350),
 .score_4 (score_4_x350),
 .score_5 (score_5_x350),
 .score_6 (score_6_x350),
 .score_7 (score_7_x350),
 .score_8 (score_8_x350),
 .score_9 (score_9_x350)
);
 
myram_28X28 #(
.ID(351),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x351),
.W_1(W_1_x351),
.W_2(W_2_x351),
.W_3(W_3_x351),
.W_4(W_4_x351),
.W_5(W_5_x351),
.W_6(W_6_x351),
.W_7(W_7_x351),
.W_8(W_8_x351),
.W_9(W_9_x351)
) u_28X28_x351 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x351),
 .score_0 (score_0_x351),
 .score_1 (score_1_x351),
 .score_2 (score_2_x351),
 .score_3 (score_3_x351),
 .score_4 (score_4_x351),
 .score_5 (score_5_x351),
 .score_6 (score_6_x351),
 .score_7 (score_7_x351),
 .score_8 (score_8_x351),
 .score_9 (score_9_x351)
);
 
myram_28X28 #(
.ID(352),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x352),
.W_1(W_1_x352),
.W_2(W_2_x352),
.W_3(W_3_x352),
.W_4(W_4_x352),
.W_5(W_5_x352),
.W_6(W_6_x352),
.W_7(W_7_x352),
.W_8(W_8_x352),
.W_9(W_9_x352)
) u_28X28_x352 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x352),
 .score_0 (score_0_x352),
 .score_1 (score_1_x352),
 .score_2 (score_2_x352),
 .score_3 (score_3_x352),
 .score_4 (score_4_x352),
 .score_5 (score_5_x352),
 .score_6 (score_6_x352),
 .score_7 (score_7_x352),
 .score_8 (score_8_x352),
 .score_9 (score_9_x352)
);
 
myram_28X28 #(
.ID(353),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x353),
.W_1(W_1_x353),
.W_2(W_2_x353),
.W_3(W_3_x353),
.W_4(W_4_x353),
.W_5(W_5_x353),
.W_6(W_6_x353),
.W_7(W_7_x353),
.W_8(W_8_x353),
.W_9(W_9_x353)
) u_28X28_x353 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x353),
 .score_0 (score_0_x353),
 .score_1 (score_1_x353),
 .score_2 (score_2_x353),
 .score_3 (score_3_x353),
 .score_4 (score_4_x353),
 .score_5 (score_5_x353),
 .score_6 (score_6_x353),
 .score_7 (score_7_x353),
 .score_8 (score_8_x353),
 .score_9 (score_9_x353)
);
 
myram_28X28 #(
.ID(354),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x354),
.W_1(W_1_x354),
.W_2(W_2_x354),
.W_3(W_3_x354),
.W_4(W_4_x354),
.W_5(W_5_x354),
.W_6(W_6_x354),
.W_7(W_7_x354),
.W_8(W_8_x354),
.W_9(W_9_x354)
) u_28X28_x354 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x354),
 .score_0 (score_0_x354),
 .score_1 (score_1_x354),
 .score_2 (score_2_x354),
 .score_3 (score_3_x354),
 .score_4 (score_4_x354),
 .score_5 (score_5_x354),
 .score_6 (score_6_x354),
 .score_7 (score_7_x354),
 .score_8 (score_8_x354),
 .score_9 (score_9_x354)
);
 
myram_28X28 #(
.ID(355),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x355),
.W_1(W_1_x355),
.W_2(W_2_x355),
.W_3(W_3_x355),
.W_4(W_4_x355),
.W_5(W_5_x355),
.W_6(W_6_x355),
.W_7(W_7_x355),
.W_8(W_8_x355),
.W_9(W_9_x355)
) u_28X28_x355 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x355),
 .score_0 (score_0_x355),
 .score_1 (score_1_x355),
 .score_2 (score_2_x355),
 .score_3 (score_3_x355),
 .score_4 (score_4_x355),
 .score_5 (score_5_x355),
 .score_6 (score_6_x355),
 .score_7 (score_7_x355),
 .score_8 (score_8_x355),
 .score_9 (score_9_x355)
);
 
myram_28X28 #(
.ID(356),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x356),
.W_1(W_1_x356),
.W_2(W_2_x356),
.W_3(W_3_x356),
.W_4(W_4_x356),
.W_5(W_5_x356),
.W_6(W_6_x356),
.W_7(W_7_x356),
.W_8(W_8_x356),
.W_9(W_9_x356)
) u_28X28_x356 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x356),
 .score_0 (score_0_x356),
 .score_1 (score_1_x356),
 .score_2 (score_2_x356),
 .score_3 (score_3_x356),
 .score_4 (score_4_x356),
 .score_5 (score_5_x356),
 .score_6 (score_6_x356),
 .score_7 (score_7_x356),
 .score_8 (score_8_x356),
 .score_9 (score_9_x356)
);
 
myram_28X28 #(
.ID(357),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x357),
.W_1(W_1_x357),
.W_2(W_2_x357),
.W_3(W_3_x357),
.W_4(W_4_x357),
.W_5(W_5_x357),
.W_6(W_6_x357),
.W_7(W_7_x357),
.W_8(W_8_x357),
.W_9(W_9_x357)
) u_28X28_x357 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x357),
 .score_0 (score_0_x357),
 .score_1 (score_1_x357),
 .score_2 (score_2_x357),
 .score_3 (score_3_x357),
 .score_4 (score_4_x357),
 .score_5 (score_5_x357),
 .score_6 (score_6_x357),
 .score_7 (score_7_x357),
 .score_8 (score_8_x357),
 .score_9 (score_9_x357)
);
 
myram_28X28 #(
.ID(358),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x358),
.W_1(W_1_x358),
.W_2(W_2_x358),
.W_3(W_3_x358),
.W_4(W_4_x358),
.W_5(W_5_x358),
.W_6(W_6_x358),
.W_7(W_7_x358),
.W_8(W_8_x358),
.W_9(W_9_x358)
) u_28X28_x358 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x358),
 .score_0 (score_0_x358),
 .score_1 (score_1_x358),
 .score_2 (score_2_x358),
 .score_3 (score_3_x358),
 .score_4 (score_4_x358),
 .score_5 (score_5_x358),
 .score_6 (score_6_x358),
 .score_7 (score_7_x358),
 .score_8 (score_8_x358),
 .score_9 (score_9_x358)
);
 
myram_28X28 #(
.ID(359),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x359),
.W_1(W_1_x359),
.W_2(W_2_x359),
.W_3(W_3_x359),
.W_4(W_4_x359),
.W_5(W_5_x359),
.W_6(W_6_x359),
.W_7(W_7_x359),
.W_8(W_8_x359),
.W_9(W_9_x359)
) u_28X28_x359 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x359),
 .score_0 (score_0_x359),
 .score_1 (score_1_x359),
 .score_2 (score_2_x359),
 .score_3 (score_3_x359),
 .score_4 (score_4_x359),
 .score_5 (score_5_x359),
 .score_6 (score_6_x359),
 .score_7 (score_7_x359),
 .score_8 (score_8_x359),
 .score_9 (score_9_x359)
);
 
myram_28X28 #(
.ID(360),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x360),
.W_1(W_1_x360),
.W_2(W_2_x360),
.W_3(W_3_x360),
.W_4(W_4_x360),
.W_5(W_5_x360),
.W_6(W_6_x360),
.W_7(W_7_x360),
.W_8(W_8_x360),
.W_9(W_9_x360)
) u_28X28_x360 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x360),
 .score_0 (score_0_x360),
 .score_1 (score_1_x360),
 .score_2 (score_2_x360),
 .score_3 (score_3_x360),
 .score_4 (score_4_x360),
 .score_5 (score_5_x360),
 .score_6 (score_6_x360),
 .score_7 (score_7_x360),
 .score_8 (score_8_x360),
 .score_9 (score_9_x360)
);
 
myram_28X28 #(
.ID(361),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x361),
.W_1(W_1_x361),
.W_2(W_2_x361),
.W_3(W_3_x361),
.W_4(W_4_x361),
.W_5(W_5_x361),
.W_6(W_6_x361),
.W_7(W_7_x361),
.W_8(W_8_x361),
.W_9(W_9_x361)
) u_28X28_x361 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x361),
 .score_0 (score_0_x361),
 .score_1 (score_1_x361),
 .score_2 (score_2_x361),
 .score_3 (score_3_x361),
 .score_4 (score_4_x361),
 .score_5 (score_5_x361),
 .score_6 (score_6_x361),
 .score_7 (score_7_x361),
 .score_8 (score_8_x361),
 .score_9 (score_9_x361)
);
 
myram_28X28 #(
.ID(362),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x362),
.W_1(W_1_x362),
.W_2(W_2_x362),
.W_3(W_3_x362),
.W_4(W_4_x362),
.W_5(W_5_x362),
.W_6(W_6_x362),
.W_7(W_7_x362),
.W_8(W_8_x362),
.W_9(W_9_x362)
) u_28X28_x362 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x362),
 .score_0 (score_0_x362),
 .score_1 (score_1_x362),
 .score_2 (score_2_x362),
 .score_3 (score_3_x362),
 .score_4 (score_4_x362),
 .score_5 (score_5_x362),
 .score_6 (score_6_x362),
 .score_7 (score_7_x362),
 .score_8 (score_8_x362),
 .score_9 (score_9_x362)
);
 
myram_28X28 #(
.ID(363),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x363),
.W_1(W_1_x363),
.W_2(W_2_x363),
.W_3(W_3_x363),
.W_4(W_4_x363),
.W_5(W_5_x363),
.W_6(W_6_x363),
.W_7(W_7_x363),
.W_8(W_8_x363),
.W_9(W_9_x363)
) u_28X28_x363 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x363),
 .score_0 (score_0_x363),
 .score_1 (score_1_x363),
 .score_2 (score_2_x363),
 .score_3 (score_3_x363),
 .score_4 (score_4_x363),
 .score_5 (score_5_x363),
 .score_6 (score_6_x363),
 .score_7 (score_7_x363),
 .score_8 (score_8_x363),
 .score_9 (score_9_x363)
);
 
myram_28X28 #(
.ID(364),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x364),
.W_1(W_1_x364),
.W_2(W_2_x364),
.W_3(W_3_x364),
.W_4(W_4_x364),
.W_5(W_5_x364),
.W_6(W_6_x364),
.W_7(W_7_x364),
.W_8(W_8_x364),
.W_9(W_9_x364)
) u_28X28_x364 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x364),
 .score_0 (score_0_x364),
 .score_1 (score_1_x364),
 .score_2 (score_2_x364),
 .score_3 (score_3_x364),
 .score_4 (score_4_x364),
 .score_5 (score_5_x364),
 .score_6 (score_6_x364),
 .score_7 (score_7_x364),
 .score_8 (score_8_x364),
 .score_9 (score_9_x364)
);
 
myram_28X28 #(
.ID(365),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x365),
.W_1(W_1_x365),
.W_2(W_2_x365),
.W_3(W_3_x365),
.W_4(W_4_x365),
.W_5(W_5_x365),
.W_6(W_6_x365),
.W_7(W_7_x365),
.W_8(W_8_x365),
.W_9(W_9_x365)
) u_28X28_x365 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x365),
 .score_0 (score_0_x365),
 .score_1 (score_1_x365),
 .score_2 (score_2_x365),
 .score_3 (score_3_x365),
 .score_4 (score_4_x365),
 .score_5 (score_5_x365),
 .score_6 (score_6_x365),
 .score_7 (score_7_x365),
 .score_8 (score_8_x365),
 .score_9 (score_9_x365)
);
 
myram_28X28 #(
.ID(366),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x366),
.W_1(W_1_x366),
.W_2(W_2_x366),
.W_3(W_3_x366),
.W_4(W_4_x366),
.W_5(W_5_x366),
.W_6(W_6_x366),
.W_7(W_7_x366),
.W_8(W_8_x366),
.W_9(W_9_x366)
) u_28X28_x366 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x366),
 .score_0 (score_0_x366),
 .score_1 (score_1_x366),
 .score_2 (score_2_x366),
 .score_3 (score_3_x366),
 .score_4 (score_4_x366),
 .score_5 (score_5_x366),
 .score_6 (score_6_x366),
 .score_7 (score_7_x366),
 .score_8 (score_8_x366),
 .score_9 (score_9_x366)
);
 
myram_28X28 #(
.ID(367),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x367),
.W_1(W_1_x367),
.W_2(W_2_x367),
.W_3(W_3_x367),
.W_4(W_4_x367),
.W_5(W_5_x367),
.W_6(W_6_x367),
.W_7(W_7_x367),
.W_8(W_8_x367),
.W_9(W_9_x367)
) u_28X28_x367 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x367),
 .score_0 (score_0_x367),
 .score_1 (score_1_x367),
 .score_2 (score_2_x367),
 .score_3 (score_3_x367),
 .score_4 (score_4_x367),
 .score_5 (score_5_x367),
 .score_6 (score_6_x367),
 .score_7 (score_7_x367),
 .score_8 (score_8_x367),
 .score_9 (score_9_x367)
);
 
myram_28X28 #(
.ID(368),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x368),
.W_1(W_1_x368),
.W_2(W_2_x368),
.W_3(W_3_x368),
.W_4(W_4_x368),
.W_5(W_5_x368),
.W_6(W_6_x368),
.W_7(W_7_x368),
.W_8(W_8_x368),
.W_9(W_9_x368)
) u_28X28_x368 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x368),
 .score_0 (score_0_x368),
 .score_1 (score_1_x368),
 .score_2 (score_2_x368),
 .score_3 (score_3_x368),
 .score_4 (score_4_x368),
 .score_5 (score_5_x368),
 .score_6 (score_6_x368),
 .score_7 (score_7_x368),
 .score_8 (score_8_x368),
 .score_9 (score_9_x368)
);
 
myram_28X28 #(
.ID(369),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x369),
.W_1(W_1_x369),
.W_2(W_2_x369),
.W_3(W_3_x369),
.W_4(W_4_x369),
.W_5(W_5_x369),
.W_6(W_6_x369),
.W_7(W_7_x369),
.W_8(W_8_x369),
.W_9(W_9_x369)
) u_28X28_x369 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x369),
 .score_0 (score_0_x369),
 .score_1 (score_1_x369),
 .score_2 (score_2_x369),
 .score_3 (score_3_x369),
 .score_4 (score_4_x369),
 .score_5 (score_5_x369),
 .score_6 (score_6_x369),
 .score_7 (score_7_x369),
 .score_8 (score_8_x369),
 .score_9 (score_9_x369)
);
 
myram_28X28 #(
.ID(370),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x370),
.W_1(W_1_x370),
.W_2(W_2_x370),
.W_3(W_3_x370),
.W_4(W_4_x370),
.W_5(W_5_x370),
.W_6(W_6_x370),
.W_7(W_7_x370),
.W_8(W_8_x370),
.W_9(W_9_x370)
) u_28X28_x370 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x370),
 .score_0 (score_0_x370),
 .score_1 (score_1_x370),
 .score_2 (score_2_x370),
 .score_3 (score_3_x370),
 .score_4 (score_4_x370),
 .score_5 (score_5_x370),
 .score_6 (score_6_x370),
 .score_7 (score_7_x370),
 .score_8 (score_8_x370),
 .score_9 (score_9_x370)
);
 
myram_28X28 #(
.ID(371),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x371),
.W_1(W_1_x371),
.W_2(W_2_x371),
.W_3(W_3_x371),
.W_4(W_4_x371),
.W_5(W_5_x371),
.W_6(W_6_x371),
.W_7(W_7_x371),
.W_8(W_8_x371),
.W_9(W_9_x371)
) u_28X28_x371 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x371),
 .score_0 (score_0_x371),
 .score_1 (score_1_x371),
 .score_2 (score_2_x371),
 .score_3 (score_3_x371),
 .score_4 (score_4_x371),
 .score_5 (score_5_x371),
 .score_6 (score_6_x371),
 .score_7 (score_7_x371),
 .score_8 (score_8_x371),
 .score_9 (score_9_x371)
);
 
myram_28X28 #(
.ID(372),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x372),
.W_1(W_1_x372),
.W_2(W_2_x372),
.W_3(W_3_x372),
.W_4(W_4_x372),
.W_5(W_5_x372),
.W_6(W_6_x372),
.W_7(W_7_x372),
.W_8(W_8_x372),
.W_9(W_9_x372)
) u_28X28_x372 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x372),
 .score_0 (score_0_x372),
 .score_1 (score_1_x372),
 .score_2 (score_2_x372),
 .score_3 (score_3_x372),
 .score_4 (score_4_x372),
 .score_5 (score_5_x372),
 .score_6 (score_6_x372),
 .score_7 (score_7_x372),
 .score_8 (score_8_x372),
 .score_9 (score_9_x372)
);
 
myram_28X28 #(
.ID(373),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x373),
.W_1(W_1_x373),
.W_2(W_2_x373),
.W_3(W_3_x373),
.W_4(W_4_x373),
.W_5(W_5_x373),
.W_6(W_6_x373),
.W_7(W_7_x373),
.W_8(W_8_x373),
.W_9(W_9_x373)
) u_28X28_x373 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x373),
 .score_0 (score_0_x373),
 .score_1 (score_1_x373),
 .score_2 (score_2_x373),
 .score_3 (score_3_x373),
 .score_4 (score_4_x373),
 .score_5 (score_5_x373),
 .score_6 (score_6_x373),
 .score_7 (score_7_x373),
 .score_8 (score_8_x373),
 .score_9 (score_9_x373)
);
 
myram_28X28 #(
.ID(374),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x374),
.W_1(W_1_x374),
.W_2(W_2_x374),
.W_3(W_3_x374),
.W_4(W_4_x374),
.W_5(W_5_x374),
.W_6(W_6_x374),
.W_7(W_7_x374),
.W_8(W_8_x374),
.W_9(W_9_x374)
) u_28X28_x374 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x374),
 .score_0 (score_0_x374),
 .score_1 (score_1_x374),
 .score_2 (score_2_x374),
 .score_3 (score_3_x374),
 .score_4 (score_4_x374),
 .score_5 (score_5_x374),
 .score_6 (score_6_x374),
 .score_7 (score_7_x374),
 .score_8 (score_8_x374),
 .score_9 (score_9_x374)
);
 
myram_28X28 #(
.ID(375),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x375),
.W_1(W_1_x375),
.W_2(W_2_x375),
.W_3(W_3_x375),
.W_4(W_4_x375),
.W_5(W_5_x375),
.W_6(W_6_x375),
.W_7(W_7_x375),
.W_8(W_8_x375),
.W_9(W_9_x375)
) u_28X28_x375 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x375),
 .score_0 (score_0_x375),
 .score_1 (score_1_x375),
 .score_2 (score_2_x375),
 .score_3 (score_3_x375),
 .score_4 (score_4_x375),
 .score_5 (score_5_x375),
 .score_6 (score_6_x375),
 .score_7 (score_7_x375),
 .score_8 (score_8_x375),
 .score_9 (score_9_x375)
);
 
myram_28X28 #(
.ID(376),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x376),
.W_1(W_1_x376),
.W_2(W_2_x376),
.W_3(W_3_x376),
.W_4(W_4_x376),
.W_5(W_5_x376),
.W_6(W_6_x376),
.W_7(W_7_x376),
.W_8(W_8_x376),
.W_9(W_9_x376)
) u_28X28_x376 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x376),
 .score_0 (score_0_x376),
 .score_1 (score_1_x376),
 .score_2 (score_2_x376),
 .score_3 (score_3_x376),
 .score_4 (score_4_x376),
 .score_5 (score_5_x376),
 .score_6 (score_6_x376),
 .score_7 (score_7_x376),
 .score_8 (score_8_x376),
 .score_9 (score_9_x376)
);
 
myram_28X28 #(
.ID(377),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x377),
.W_1(W_1_x377),
.W_2(W_2_x377),
.W_3(W_3_x377),
.W_4(W_4_x377),
.W_5(W_5_x377),
.W_6(W_6_x377),
.W_7(W_7_x377),
.W_8(W_8_x377),
.W_9(W_9_x377)
) u_28X28_x377 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x377),
 .score_0 (score_0_x377),
 .score_1 (score_1_x377),
 .score_2 (score_2_x377),
 .score_3 (score_3_x377),
 .score_4 (score_4_x377),
 .score_5 (score_5_x377),
 .score_6 (score_6_x377),
 .score_7 (score_7_x377),
 .score_8 (score_8_x377),
 .score_9 (score_9_x377)
);
 
myram_28X28 #(
.ID(378),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x378),
.W_1(W_1_x378),
.W_2(W_2_x378),
.W_3(W_3_x378),
.W_4(W_4_x378),
.W_5(W_5_x378),
.W_6(W_6_x378),
.W_7(W_7_x378),
.W_8(W_8_x378),
.W_9(W_9_x378)
) u_28X28_x378 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x378),
 .score_0 (score_0_x378),
 .score_1 (score_1_x378),
 .score_2 (score_2_x378),
 .score_3 (score_3_x378),
 .score_4 (score_4_x378),
 .score_5 (score_5_x378),
 .score_6 (score_6_x378),
 .score_7 (score_7_x378),
 .score_8 (score_8_x378),
 .score_9 (score_9_x378)
);
 
myram_28X28 #(
.ID(379),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x379),
.W_1(W_1_x379),
.W_2(W_2_x379),
.W_3(W_3_x379),
.W_4(W_4_x379),
.W_5(W_5_x379),
.W_6(W_6_x379),
.W_7(W_7_x379),
.W_8(W_8_x379),
.W_9(W_9_x379)
) u_28X28_x379 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x379),
 .score_0 (score_0_x379),
 .score_1 (score_1_x379),
 .score_2 (score_2_x379),
 .score_3 (score_3_x379),
 .score_4 (score_4_x379),
 .score_5 (score_5_x379),
 .score_6 (score_6_x379),
 .score_7 (score_7_x379),
 .score_8 (score_8_x379),
 .score_9 (score_9_x379)
);
 
myram_28X28 #(
.ID(380),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x380),
.W_1(W_1_x380),
.W_2(W_2_x380),
.W_3(W_3_x380),
.W_4(W_4_x380),
.W_5(W_5_x380),
.W_6(W_6_x380),
.W_7(W_7_x380),
.W_8(W_8_x380),
.W_9(W_9_x380)
) u_28X28_x380 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x380),
 .score_0 (score_0_x380),
 .score_1 (score_1_x380),
 .score_2 (score_2_x380),
 .score_3 (score_3_x380),
 .score_4 (score_4_x380),
 .score_5 (score_5_x380),
 .score_6 (score_6_x380),
 .score_7 (score_7_x380),
 .score_8 (score_8_x380),
 .score_9 (score_9_x380)
);
 
myram_28X28 #(
.ID(381),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x381),
.W_1(W_1_x381),
.W_2(W_2_x381),
.W_3(W_3_x381),
.W_4(W_4_x381),
.W_5(W_5_x381),
.W_6(W_6_x381),
.W_7(W_7_x381),
.W_8(W_8_x381),
.W_9(W_9_x381)
) u_28X28_x381 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x381),
 .score_0 (score_0_x381),
 .score_1 (score_1_x381),
 .score_2 (score_2_x381),
 .score_3 (score_3_x381),
 .score_4 (score_4_x381),
 .score_5 (score_5_x381),
 .score_6 (score_6_x381),
 .score_7 (score_7_x381),
 .score_8 (score_8_x381),
 .score_9 (score_9_x381)
);
 
myram_28X28 #(
.ID(382),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x382),
.W_1(W_1_x382),
.W_2(W_2_x382),
.W_3(W_3_x382),
.W_4(W_4_x382),
.W_5(W_5_x382),
.W_6(W_6_x382),
.W_7(W_7_x382),
.W_8(W_8_x382),
.W_9(W_9_x382)
) u_28X28_x382 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x382),
 .score_0 (score_0_x382),
 .score_1 (score_1_x382),
 .score_2 (score_2_x382),
 .score_3 (score_3_x382),
 .score_4 (score_4_x382),
 .score_5 (score_5_x382),
 .score_6 (score_6_x382),
 .score_7 (score_7_x382),
 .score_8 (score_8_x382),
 .score_9 (score_9_x382)
);
 
myram_28X28 #(
.ID(383),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x383),
.W_1(W_1_x383),
.W_2(W_2_x383),
.W_3(W_3_x383),
.W_4(W_4_x383),
.W_5(W_5_x383),
.W_6(W_6_x383),
.W_7(W_7_x383),
.W_8(W_8_x383),
.W_9(W_9_x383)
) u_28X28_x383 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x383),
 .score_0 (score_0_x383),
 .score_1 (score_1_x383),
 .score_2 (score_2_x383),
 .score_3 (score_3_x383),
 .score_4 (score_4_x383),
 .score_5 (score_5_x383),
 .score_6 (score_6_x383),
 .score_7 (score_7_x383),
 .score_8 (score_8_x383),
 .score_9 (score_9_x383)
);
 
myram_28X28 #(
.ID(384),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x384),
.W_1(W_1_x384),
.W_2(W_2_x384),
.W_3(W_3_x384),
.W_4(W_4_x384),
.W_5(W_5_x384),
.W_6(W_6_x384),
.W_7(W_7_x384),
.W_8(W_8_x384),
.W_9(W_9_x384)
) u_28X28_x384 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x384),
 .score_0 (score_0_x384),
 .score_1 (score_1_x384),
 .score_2 (score_2_x384),
 .score_3 (score_3_x384),
 .score_4 (score_4_x384),
 .score_5 (score_5_x384),
 .score_6 (score_6_x384),
 .score_7 (score_7_x384),
 .score_8 (score_8_x384),
 .score_9 (score_9_x384)
);
 
myram_28X28 #(
.ID(385),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x385),
.W_1(W_1_x385),
.W_2(W_2_x385),
.W_3(W_3_x385),
.W_4(W_4_x385),
.W_5(W_5_x385),
.W_6(W_6_x385),
.W_7(W_7_x385),
.W_8(W_8_x385),
.W_9(W_9_x385)
) u_28X28_x385 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x385),
 .score_0 (score_0_x385),
 .score_1 (score_1_x385),
 .score_2 (score_2_x385),
 .score_3 (score_3_x385),
 .score_4 (score_4_x385),
 .score_5 (score_5_x385),
 .score_6 (score_6_x385),
 .score_7 (score_7_x385),
 .score_8 (score_8_x385),
 .score_9 (score_9_x385)
);
 
myram_28X28 #(
.ID(386),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x386),
.W_1(W_1_x386),
.W_2(W_2_x386),
.W_3(W_3_x386),
.W_4(W_4_x386),
.W_5(W_5_x386),
.W_6(W_6_x386),
.W_7(W_7_x386),
.W_8(W_8_x386),
.W_9(W_9_x386)
) u_28X28_x386 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x386),
 .score_0 (score_0_x386),
 .score_1 (score_1_x386),
 .score_2 (score_2_x386),
 .score_3 (score_3_x386),
 .score_4 (score_4_x386),
 .score_5 (score_5_x386),
 .score_6 (score_6_x386),
 .score_7 (score_7_x386),
 .score_8 (score_8_x386),
 .score_9 (score_9_x386)
);
 
myram_28X28 #(
.ID(387),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x387),
.W_1(W_1_x387),
.W_2(W_2_x387),
.W_3(W_3_x387),
.W_4(W_4_x387),
.W_5(W_5_x387),
.W_6(W_6_x387),
.W_7(W_7_x387),
.W_8(W_8_x387),
.W_9(W_9_x387)
) u_28X28_x387 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x387),
 .score_0 (score_0_x387),
 .score_1 (score_1_x387),
 .score_2 (score_2_x387),
 .score_3 (score_3_x387),
 .score_4 (score_4_x387),
 .score_5 (score_5_x387),
 .score_6 (score_6_x387),
 .score_7 (score_7_x387),
 .score_8 (score_8_x387),
 .score_9 (score_9_x387)
);
 
myram_28X28 #(
.ID(388),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x388),
.W_1(W_1_x388),
.W_2(W_2_x388),
.W_3(W_3_x388),
.W_4(W_4_x388),
.W_5(W_5_x388),
.W_6(W_6_x388),
.W_7(W_7_x388),
.W_8(W_8_x388),
.W_9(W_9_x388)
) u_28X28_x388 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x388),
 .score_0 (score_0_x388),
 .score_1 (score_1_x388),
 .score_2 (score_2_x388),
 .score_3 (score_3_x388),
 .score_4 (score_4_x388),
 .score_5 (score_5_x388),
 .score_6 (score_6_x388),
 .score_7 (score_7_x388),
 .score_8 (score_8_x388),
 .score_9 (score_9_x388)
);
 
myram_28X28 #(
.ID(389),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x389),
.W_1(W_1_x389),
.W_2(W_2_x389),
.W_3(W_3_x389),
.W_4(W_4_x389),
.W_5(W_5_x389),
.W_6(W_6_x389),
.W_7(W_7_x389),
.W_8(W_8_x389),
.W_9(W_9_x389)
) u_28X28_x389 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x389),
 .score_0 (score_0_x389),
 .score_1 (score_1_x389),
 .score_2 (score_2_x389),
 .score_3 (score_3_x389),
 .score_4 (score_4_x389),
 .score_5 (score_5_x389),
 .score_6 (score_6_x389),
 .score_7 (score_7_x389),
 .score_8 (score_8_x389),
 .score_9 (score_9_x389)
);
 
myram_28X28 #(
.ID(390),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x390),
.W_1(W_1_x390),
.W_2(W_2_x390),
.W_3(W_3_x390),
.W_4(W_4_x390),
.W_5(W_5_x390),
.W_6(W_6_x390),
.W_7(W_7_x390),
.W_8(W_8_x390),
.W_9(W_9_x390)
) u_28X28_x390 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x390),
 .score_0 (score_0_x390),
 .score_1 (score_1_x390),
 .score_2 (score_2_x390),
 .score_3 (score_3_x390),
 .score_4 (score_4_x390),
 .score_5 (score_5_x390),
 .score_6 (score_6_x390),
 .score_7 (score_7_x390),
 .score_8 (score_8_x390),
 .score_9 (score_9_x390)
);
 
myram_28X28 #(
.ID(391),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x391),
.W_1(W_1_x391),
.W_2(W_2_x391),
.W_3(W_3_x391),
.W_4(W_4_x391),
.W_5(W_5_x391),
.W_6(W_6_x391),
.W_7(W_7_x391),
.W_8(W_8_x391),
.W_9(W_9_x391)
) u_28X28_x391 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x391),
 .score_0 (score_0_x391),
 .score_1 (score_1_x391),
 .score_2 (score_2_x391),
 .score_3 (score_3_x391),
 .score_4 (score_4_x391),
 .score_5 (score_5_x391),
 .score_6 (score_6_x391),
 .score_7 (score_7_x391),
 .score_8 (score_8_x391),
 .score_9 (score_9_x391)
);
 
myram_28X28 #(
.ID(392),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x392),
.W_1(W_1_x392),
.W_2(W_2_x392),
.W_3(W_3_x392),
.W_4(W_4_x392),
.W_5(W_5_x392),
.W_6(W_6_x392),
.W_7(W_7_x392),
.W_8(W_8_x392),
.W_9(W_9_x392)
) u_28X28_x392 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x392),
 .score_0 (score_0_x392),
 .score_1 (score_1_x392),
 .score_2 (score_2_x392),
 .score_3 (score_3_x392),
 .score_4 (score_4_x392),
 .score_5 (score_5_x392),
 .score_6 (score_6_x392),
 .score_7 (score_7_x392),
 .score_8 (score_8_x392),
 .score_9 (score_9_x392)
);
 
myram_28X28 #(
.ID(393),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x393),
.W_1(W_1_x393),
.W_2(W_2_x393),
.W_3(W_3_x393),
.W_4(W_4_x393),
.W_5(W_5_x393),
.W_6(W_6_x393),
.W_7(W_7_x393),
.W_8(W_8_x393),
.W_9(W_9_x393)
) u_28X28_x393 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x393),
 .score_0 (score_0_x393),
 .score_1 (score_1_x393),
 .score_2 (score_2_x393),
 .score_3 (score_3_x393),
 .score_4 (score_4_x393),
 .score_5 (score_5_x393),
 .score_6 (score_6_x393),
 .score_7 (score_7_x393),
 .score_8 (score_8_x393),
 .score_9 (score_9_x393)
);
 
myram_28X28 #(
.ID(394),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x394),
.W_1(W_1_x394),
.W_2(W_2_x394),
.W_3(W_3_x394),
.W_4(W_4_x394),
.W_5(W_5_x394),
.W_6(W_6_x394),
.W_7(W_7_x394),
.W_8(W_8_x394),
.W_9(W_9_x394)
) u_28X28_x394 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x394),
 .score_0 (score_0_x394),
 .score_1 (score_1_x394),
 .score_2 (score_2_x394),
 .score_3 (score_3_x394),
 .score_4 (score_4_x394),
 .score_5 (score_5_x394),
 .score_6 (score_6_x394),
 .score_7 (score_7_x394),
 .score_8 (score_8_x394),
 .score_9 (score_9_x394)
);
 
myram_28X28 #(
.ID(395),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x395),
.W_1(W_1_x395),
.W_2(W_2_x395),
.W_3(W_3_x395),
.W_4(W_4_x395),
.W_5(W_5_x395),
.W_6(W_6_x395),
.W_7(W_7_x395),
.W_8(W_8_x395),
.W_9(W_9_x395)
) u_28X28_x395 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x395),
 .score_0 (score_0_x395),
 .score_1 (score_1_x395),
 .score_2 (score_2_x395),
 .score_3 (score_3_x395),
 .score_4 (score_4_x395),
 .score_5 (score_5_x395),
 .score_6 (score_6_x395),
 .score_7 (score_7_x395),
 .score_8 (score_8_x395),
 .score_9 (score_9_x395)
);
 
myram_28X28 #(
.ID(396),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x396),
.W_1(W_1_x396),
.W_2(W_2_x396),
.W_3(W_3_x396),
.W_4(W_4_x396),
.W_5(W_5_x396),
.W_6(W_6_x396),
.W_7(W_7_x396),
.W_8(W_8_x396),
.W_9(W_9_x396)
) u_28X28_x396 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x396),
 .score_0 (score_0_x396),
 .score_1 (score_1_x396),
 .score_2 (score_2_x396),
 .score_3 (score_3_x396),
 .score_4 (score_4_x396),
 .score_5 (score_5_x396),
 .score_6 (score_6_x396),
 .score_7 (score_7_x396),
 .score_8 (score_8_x396),
 .score_9 (score_9_x396)
);
 
myram_28X28 #(
.ID(397),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x397),
.W_1(W_1_x397),
.W_2(W_2_x397),
.W_3(W_3_x397),
.W_4(W_4_x397),
.W_5(W_5_x397),
.W_6(W_6_x397),
.W_7(W_7_x397),
.W_8(W_8_x397),
.W_9(W_9_x397)
) u_28X28_x397 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x397),
 .score_0 (score_0_x397),
 .score_1 (score_1_x397),
 .score_2 (score_2_x397),
 .score_3 (score_3_x397),
 .score_4 (score_4_x397),
 .score_5 (score_5_x397),
 .score_6 (score_6_x397),
 .score_7 (score_7_x397),
 .score_8 (score_8_x397),
 .score_9 (score_9_x397)
);
 
myram_28X28 #(
.ID(398),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x398),
.W_1(W_1_x398),
.W_2(W_2_x398),
.W_3(W_3_x398),
.W_4(W_4_x398),
.W_5(W_5_x398),
.W_6(W_6_x398),
.W_7(W_7_x398),
.W_8(W_8_x398),
.W_9(W_9_x398)
) u_28X28_x398 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x398),
 .score_0 (score_0_x398),
 .score_1 (score_1_x398),
 .score_2 (score_2_x398),
 .score_3 (score_3_x398),
 .score_4 (score_4_x398),
 .score_5 (score_5_x398),
 .score_6 (score_6_x398),
 .score_7 (score_7_x398),
 .score_8 (score_8_x398),
 .score_9 (score_9_x398)
);
 
myram_28X28 #(
.ID(399),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x399),
.W_1(W_1_x399),
.W_2(W_2_x399),
.W_3(W_3_x399),
.W_4(W_4_x399),
.W_5(W_5_x399),
.W_6(W_6_x399),
.W_7(W_7_x399),
.W_8(W_8_x399),
.W_9(W_9_x399)
) u_28X28_x399 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x399),
 .score_0 (score_0_x399),
 .score_1 (score_1_x399),
 .score_2 (score_2_x399),
 .score_3 (score_3_x399),
 .score_4 (score_4_x399),
 .score_5 (score_5_x399),
 .score_6 (score_6_x399),
 .score_7 (score_7_x399),
 .score_8 (score_8_x399),
 .score_9 (score_9_x399)
);
 
myram_28X28 #(
.ID(400),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x400),
.W_1(W_1_x400),
.W_2(W_2_x400),
.W_3(W_3_x400),
.W_4(W_4_x400),
.W_5(W_5_x400),
.W_6(W_6_x400),
.W_7(W_7_x400),
.W_8(W_8_x400),
.W_9(W_9_x400)
) u_28X28_x400 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x400),
 .score_0 (score_0_x400),
 .score_1 (score_1_x400),
 .score_2 (score_2_x400),
 .score_3 (score_3_x400),
 .score_4 (score_4_x400),
 .score_5 (score_5_x400),
 .score_6 (score_6_x400),
 .score_7 (score_7_x400),
 .score_8 (score_8_x400),
 .score_9 (score_9_x400)
);
 
myram_28X28 #(
.ID(401),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x401),
.W_1(W_1_x401),
.W_2(W_2_x401),
.W_3(W_3_x401),
.W_4(W_4_x401),
.W_5(W_5_x401),
.W_6(W_6_x401),
.W_7(W_7_x401),
.W_8(W_8_x401),
.W_9(W_9_x401)
) u_28X28_x401 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x401),
 .score_0 (score_0_x401),
 .score_1 (score_1_x401),
 .score_2 (score_2_x401),
 .score_3 (score_3_x401),
 .score_4 (score_4_x401),
 .score_5 (score_5_x401),
 .score_6 (score_6_x401),
 .score_7 (score_7_x401),
 .score_8 (score_8_x401),
 .score_9 (score_9_x401)
);
 
myram_28X28 #(
.ID(402),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x402),
.W_1(W_1_x402),
.W_2(W_2_x402),
.W_3(W_3_x402),
.W_4(W_4_x402),
.W_5(W_5_x402),
.W_6(W_6_x402),
.W_7(W_7_x402),
.W_8(W_8_x402),
.W_9(W_9_x402)
) u_28X28_x402 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x402),
 .score_0 (score_0_x402),
 .score_1 (score_1_x402),
 .score_2 (score_2_x402),
 .score_3 (score_3_x402),
 .score_4 (score_4_x402),
 .score_5 (score_5_x402),
 .score_6 (score_6_x402),
 .score_7 (score_7_x402),
 .score_8 (score_8_x402),
 .score_9 (score_9_x402)
);
 
myram_28X28 #(
.ID(403),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x403),
.W_1(W_1_x403),
.W_2(W_2_x403),
.W_3(W_3_x403),
.W_4(W_4_x403),
.W_5(W_5_x403),
.W_6(W_6_x403),
.W_7(W_7_x403),
.W_8(W_8_x403),
.W_9(W_9_x403)
) u_28X28_x403 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x403),
 .score_0 (score_0_x403),
 .score_1 (score_1_x403),
 .score_2 (score_2_x403),
 .score_3 (score_3_x403),
 .score_4 (score_4_x403),
 .score_5 (score_5_x403),
 .score_6 (score_6_x403),
 .score_7 (score_7_x403),
 .score_8 (score_8_x403),
 .score_9 (score_9_x403)
);
 
myram_28X28 #(
.ID(404),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x404),
.W_1(W_1_x404),
.W_2(W_2_x404),
.W_3(W_3_x404),
.W_4(W_4_x404),
.W_5(W_5_x404),
.W_6(W_6_x404),
.W_7(W_7_x404),
.W_8(W_8_x404),
.W_9(W_9_x404)
) u_28X28_x404 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x404),
 .score_0 (score_0_x404),
 .score_1 (score_1_x404),
 .score_2 (score_2_x404),
 .score_3 (score_3_x404),
 .score_4 (score_4_x404),
 .score_5 (score_5_x404),
 .score_6 (score_6_x404),
 .score_7 (score_7_x404),
 .score_8 (score_8_x404),
 .score_9 (score_9_x404)
);
 
myram_28X28 #(
.ID(405),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x405),
.W_1(W_1_x405),
.W_2(W_2_x405),
.W_3(W_3_x405),
.W_4(W_4_x405),
.W_5(W_5_x405),
.W_6(W_6_x405),
.W_7(W_7_x405),
.W_8(W_8_x405),
.W_9(W_9_x405)
) u_28X28_x405 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x405),
 .score_0 (score_0_x405),
 .score_1 (score_1_x405),
 .score_2 (score_2_x405),
 .score_3 (score_3_x405),
 .score_4 (score_4_x405),
 .score_5 (score_5_x405),
 .score_6 (score_6_x405),
 .score_7 (score_7_x405),
 .score_8 (score_8_x405),
 .score_9 (score_9_x405)
);
 
myram_28X28 #(
.ID(406),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x406),
.W_1(W_1_x406),
.W_2(W_2_x406),
.W_3(W_3_x406),
.W_4(W_4_x406),
.W_5(W_5_x406),
.W_6(W_6_x406),
.W_7(W_7_x406),
.W_8(W_8_x406),
.W_9(W_9_x406)
) u_28X28_x406 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x406),
 .score_0 (score_0_x406),
 .score_1 (score_1_x406),
 .score_2 (score_2_x406),
 .score_3 (score_3_x406),
 .score_4 (score_4_x406),
 .score_5 (score_5_x406),
 .score_6 (score_6_x406),
 .score_7 (score_7_x406),
 .score_8 (score_8_x406),
 .score_9 (score_9_x406)
);
 
myram_28X28 #(
.ID(407),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x407),
.W_1(W_1_x407),
.W_2(W_2_x407),
.W_3(W_3_x407),
.W_4(W_4_x407),
.W_5(W_5_x407),
.W_6(W_6_x407),
.W_7(W_7_x407),
.W_8(W_8_x407),
.W_9(W_9_x407)
) u_28X28_x407 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x407),
 .score_0 (score_0_x407),
 .score_1 (score_1_x407),
 .score_2 (score_2_x407),
 .score_3 (score_3_x407),
 .score_4 (score_4_x407),
 .score_5 (score_5_x407),
 .score_6 (score_6_x407),
 .score_7 (score_7_x407),
 .score_8 (score_8_x407),
 .score_9 (score_9_x407)
);
 
myram_28X28 #(
.ID(408),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x408),
.W_1(W_1_x408),
.W_2(W_2_x408),
.W_3(W_3_x408),
.W_4(W_4_x408),
.W_5(W_5_x408),
.W_6(W_6_x408),
.W_7(W_7_x408),
.W_8(W_8_x408),
.W_9(W_9_x408)
) u_28X28_x408 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x408),
 .score_0 (score_0_x408),
 .score_1 (score_1_x408),
 .score_2 (score_2_x408),
 .score_3 (score_3_x408),
 .score_4 (score_4_x408),
 .score_5 (score_5_x408),
 .score_6 (score_6_x408),
 .score_7 (score_7_x408),
 .score_8 (score_8_x408),
 .score_9 (score_9_x408)
);
 
myram_28X28 #(
.ID(409),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x409),
.W_1(W_1_x409),
.W_2(W_2_x409),
.W_3(W_3_x409),
.W_4(W_4_x409),
.W_5(W_5_x409),
.W_6(W_6_x409),
.W_7(W_7_x409),
.W_8(W_8_x409),
.W_9(W_9_x409)
) u_28X28_x409 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x409),
 .score_0 (score_0_x409),
 .score_1 (score_1_x409),
 .score_2 (score_2_x409),
 .score_3 (score_3_x409),
 .score_4 (score_4_x409),
 .score_5 (score_5_x409),
 .score_6 (score_6_x409),
 .score_7 (score_7_x409),
 .score_8 (score_8_x409),
 .score_9 (score_9_x409)
);
 
myram_28X28 #(
.ID(410),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x410),
.W_1(W_1_x410),
.W_2(W_2_x410),
.W_3(W_3_x410),
.W_4(W_4_x410),
.W_5(W_5_x410),
.W_6(W_6_x410),
.W_7(W_7_x410),
.W_8(W_8_x410),
.W_9(W_9_x410)
) u_28X28_x410 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x410),
 .score_0 (score_0_x410),
 .score_1 (score_1_x410),
 .score_2 (score_2_x410),
 .score_3 (score_3_x410),
 .score_4 (score_4_x410),
 .score_5 (score_5_x410),
 .score_6 (score_6_x410),
 .score_7 (score_7_x410),
 .score_8 (score_8_x410),
 .score_9 (score_9_x410)
);
 
myram_28X28 #(
.ID(411),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x411),
.W_1(W_1_x411),
.W_2(W_2_x411),
.W_3(W_3_x411),
.W_4(W_4_x411),
.W_5(W_5_x411),
.W_6(W_6_x411),
.W_7(W_7_x411),
.W_8(W_8_x411),
.W_9(W_9_x411)
) u_28X28_x411 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x411),
 .score_0 (score_0_x411),
 .score_1 (score_1_x411),
 .score_2 (score_2_x411),
 .score_3 (score_3_x411),
 .score_4 (score_4_x411),
 .score_5 (score_5_x411),
 .score_6 (score_6_x411),
 .score_7 (score_7_x411),
 .score_8 (score_8_x411),
 .score_9 (score_9_x411)
);
 
myram_28X28 #(
.ID(412),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x412),
.W_1(W_1_x412),
.W_2(W_2_x412),
.W_3(W_3_x412),
.W_4(W_4_x412),
.W_5(W_5_x412),
.W_6(W_6_x412),
.W_7(W_7_x412),
.W_8(W_8_x412),
.W_9(W_9_x412)
) u_28X28_x412 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x412),
 .score_0 (score_0_x412),
 .score_1 (score_1_x412),
 .score_2 (score_2_x412),
 .score_3 (score_3_x412),
 .score_4 (score_4_x412),
 .score_5 (score_5_x412),
 .score_6 (score_6_x412),
 .score_7 (score_7_x412),
 .score_8 (score_8_x412),
 .score_9 (score_9_x412)
);
 
myram_28X28 #(
.ID(413),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x413),
.W_1(W_1_x413),
.W_2(W_2_x413),
.W_3(W_3_x413),
.W_4(W_4_x413),
.W_5(W_5_x413),
.W_6(W_6_x413),
.W_7(W_7_x413),
.W_8(W_8_x413),
.W_9(W_9_x413)
) u_28X28_x413 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x413),
 .score_0 (score_0_x413),
 .score_1 (score_1_x413),
 .score_2 (score_2_x413),
 .score_3 (score_3_x413),
 .score_4 (score_4_x413),
 .score_5 (score_5_x413),
 .score_6 (score_6_x413),
 .score_7 (score_7_x413),
 .score_8 (score_8_x413),
 .score_9 (score_9_x413)
);
 
myram_28X28 #(
.ID(414),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x414),
.W_1(W_1_x414),
.W_2(W_2_x414),
.W_3(W_3_x414),
.W_4(W_4_x414),
.W_5(W_5_x414),
.W_6(W_6_x414),
.W_7(W_7_x414),
.W_8(W_8_x414),
.W_9(W_9_x414)
) u_28X28_x414 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x414),
 .score_0 (score_0_x414),
 .score_1 (score_1_x414),
 .score_2 (score_2_x414),
 .score_3 (score_3_x414),
 .score_4 (score_4_x414),
 .score_5 (score_5_x414),
 .score_6 (score_6_x414),
 .score_7 (score_7_x414),
 .score_8 (score_8_x414),
 .score_9 (score_9_x414)
);
 
myram_28X28 #(
.ID(415),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x415),
.W_1(W_1_x415),
.W_2(W_2_x415),
.W_3(W_3_x415),
.W_4(W_4_x415),
.W_5(W_5_x415),
.W_6(W_6_x415),
.W_7(W_7_x415),
.W_8(W_8_x415),
.W_9(W_9_x415)
) u_28X28_x415 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x415),
 .score_0 (score_0_x415),
 .score_1 (score_1_x415),
 .score_2 (score_2_x415),
 .score_3 (score_3_x415),
 .score_4 (score_4_x415),
 .score_5 (score_5_x415),
 .score_6 (score_6_x415),
 .score_7 (score_7_x415),
 .score_8 (score_8_x415),
 .score_9 (score_9_x415)
);
 
myram_28X28 #(
.ID(416),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x416),
.W_1(W_1_x416),
.W_2(W_2_x416),
.W_3(W_3_x416),
.W_4(W_4_x416),
.W_5(W_5_x416),
.W_6(W_6_x416),
.W_7(W_7_x416),
.W_8(W_8_x416),
.W_9(W_9_x416)
) u_28X28_x416 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x416),
 .score_0 (score_0_x416),
 .score_1 (score_1_x416),
 .score_2 (score_2_x416),
 .score_3 (score_3_x416),
 .score_4 (score_4_x416),
 .score_5 (score_5_x416),
 .score_6 (score_6_x416),
 .score_7 (score_7_x416),
 .score_8 (score_8_x416),
 .score_9 (score_9_x416)
);
 
myram_28X28 #(
.ID(417),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x417),
.W_1(W_1_x417),
.W_2(W_2_x417),
.W_3(W_3_x417),
.W_4(W_4_x417),
.W_5(W_5_x417),
.W_6(W_6_x417),
.W_7(W_7_x417),
.W_8(W_8_x417),
.W_9(W_9_x417)
) u_28X28_x417 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x417),
 .score_0 (score_0_x417),
 .score_1 (score_1_x417),
 .score_2 (score_2_x417),
 .score_3 (score_3_x417),
 .score_4 (score_4_x417),
 .score_5 (score_5_x417),
 .score_6 (score_6_x417),
 .score_7 (score_7_x417),
 .score_8 (score_8_x417),
 .score_9 (score_9_x417)
);
 
myram_28X28 #(
.ID(418),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x418),
.W_1(W_1_x418),
.W_2(W_2_x418),
.W_3(W_3_x418),
.W_4(W_4_x418),
.W_5(W_5_x418),
.W_6(W_6_x418),
.W_7(W_7_x418),
.W_8(W_8_x418),
.W_9(W_9_x418)
) u_28X28_x418 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x418),
 .score_0 (score_0_x418),
 .score_1 (score_1_x418),
 .score_2 (score_2_x418),
 .score_3 (score_3_x418),
 .score_4 (score_4_x418),
 .score_5 (score_5_x418),
 .score_6 (score_6_x418),
 .score_7 (score_7_x418),
 .score_8 (score_8_x418),
 .score_9 (score_9_x418)
);
 
myram_28X28 #(
.ID(419),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x419),
.W_1(W_1_x419),
.W_2(W_2_x419),
.W_3(W_3_x419),
.W_4(W_4_x419),
.W_5(W_5_x419),
.W_6(W_6_x419),
.W_7(W_7_x419),
.W_8(W_8_x419),
.W_9(W_9_x419)
) u_28X28_x419 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x419),
 .score_0 (score_0_x419),
 .score_1 (score_1_x419),
 .score_2 (score_2_x419),
 .score_3 (score_3_x419),
 .score_4 (score_4_x419),
 .score_5 (score_5_x419),
 .score_6 (score_6_x419),
 .score_7 (score_7_x419),
 .score_8 (score_8_x419),
 .score_9 (score_9_x419)
);
 
myram_28X28 #(
.ID(420),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x420),
.W_1(W_1_x420),
.W_2(W_2_x420),
.W_3(W_3_x420),
.W_4(W_4_x420),
.W_5(W_5_x420),
.W_6(W_6_x420),
.W_7(W_7_x420),
.W_8(W_8_x420),
.W_9(W_9_x420)
) u_28X28_x420 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x420),
 .score_0 (score_0_x420),
 .score_1 (score_1_x420),
 .score_2 (score_2_x420),
 .score_3 (score_3_x420),
 .score_4 (score_4_x420),
 .score_5 (score_5_x420),
 .score_6 (score_6_x420),
 .score_7 (score_7_x420),
 .score_8 (score_8_x420),
 .score_9 (score_9_x420)
);
 
myram_28X28 #(
.ID(421),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x421),
.W_1(W_1_x421),
.W_2(W_2_x421),
.W_3(W_3_x421),
.W_4(W_4_x421),
.W_5(W_5_x421),
.W_6(W_6_x421),
.W_7(W_7_x421),
.W_8(W_8_x421),
.W_9(W_9_x421)
) u_28X28_x421 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x421),
 .score_0 (score_0_x421),
 .score_1 (score_1_x421),
 .score_2 (score_2_x421),
 .score_3 (score_3_x421),
 .score_4 (score_4_x421),
 .score_5 (score_5_x421),
 .score_6 (score_6_x421),
 .score_7 (score_7_x421),
 .score_8 (score_8_x421),
 .score_9 (score_9_x421)
);
 
myram_28X28 #(
.ID(422),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x422),
.W_1(W_1_x422),
.W_2(W_2_x422),
.W_3(W_3_x422),
.W_4(W_4_x422),
.W_5(W_5_x422),
.W_6(W_6_x422),
.W_7(W_7_x422),
.W_8(W_8_x422),
.W_9(W_9_x422)
) u_28X28_x422 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x422),
 .score_0 (score_0_x422),
 .score_1 (score_1_x422),
 .score_2 (score_2_x422),
 .score_3 (score_3_x422),
 .score_4 (score_4_x422),
 .score_5 (score_5_x422),
 .score_6 (score_6_x422),
 .score_7 (score_7_x422),
 .score_8 (score_8_x422),
 .score_9 (score_9_x422)
);
 
myram_28X28 #(
.ID(423),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x423),
.W_1(W_1_x423),
.W_2(W_2_x423),
.W_3(W_3_x423),
.W_4(W_4_x423),
.W_5(W_5_x423),
.W_6(W_6_x423),
.W_7(W_7_x423),
.W_8(W_8_x423),
.W_9(W_9_x423)
) u_28X28_x423 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x423),
 .score_0 (score_0_x423),
 .score_1 (score_1_x423),
 .score_2 (score_2_x423),
 .score_3 (score_3_x423),
 .score_4 (score_4_x423),
 .score_5 (score_5_x423),
 .score_6 (score_6_x423),
 .score_7 (score_7_x423),
 .score_8 (score_8_x423),
 .score_9 (score_9_x423)
);
 
myram_28X28 #(
.ID(424),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x424),
.W_1(W_1_x424),
.W_2(W_2_x424),
.W_3(W_3_x424),
.W_4(W_4_x424),
.W_5(W_5_x424),
.W_6(W_6_x424),
.W_7(W_7_x424),
.W_8(W_8_x424),
.W_9(W_9_x424)
) u_28X28_x424 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x424),
 .score_0 (score_0_x424),
 .score_1 (score_1_x424),
 .score_2 (score_2_x424),
 .score_3 (score_3_x424),
 .score_4 (score_4_x424),
 .score_5 (score_5_x424),
 .score_6 (score_6_x424),
 .score_7 (score_7_x424),
 .score_8 (score_8_x424),
 .score_9 (score_9_x424)
);
 
myram_28X28 #(
.ID(425),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x425),
.W_1(W_1_x425),
.W_2(W_2_x425),
.W_3(W_3_x425),
.W_4(W_4_x425),
.W_5(W_5_x425),
.W_6(W_6_x425),
.W_7(W_7_x425),
.W_8(W_8_x425),
.W_9(W_9_x425)
) u_28X28_x425 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x425),
 .score_0 (score_0_x425),
 .score_1 (score_1_x425),
 .score_2 (score_2_x425),
 .score_3 (score_3_x425),
 .score_4 (score_4_x425),
 .score_5 (score_5_x425),
 .score_6 (score_6_x425),
 .score_7 (score_7_x425),
 .score_8 (score_8_x425),
 .score_9 (score_9_x425)
);
 
myram_28X28 #(
.ID(426),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x426),
.W_1(W_1_x426),
.W_2(W_2_x426),
.W_3(W_3_x426),
.W_4(W_4_x426),
.W_5(W_5_x426),
.W_6(W_6_x426),
.W_7(W_7_x426),
.W_8(W_8_x426),
.W_9(W_9_x426)
) u_28X28_x426 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x426),
 .score_0 (score_0_x426),
 .score_1 (score_1_x426),
 .score_2 (score_2_x426),
 .score_3 (score_3_x426),
 .score_4 (score_4_x426),
 .score_5 (score_5_x426),
 .score_6 (score_6_x426),
 .score_7 (score_7_x426),
 .score_8 (score_8_x426),
 .score_9 (score_9_x426)
);
 
myram_28X28 #(
.ID(427),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x427),
.W_1(W_1_x427),
.W_2(W_2_x427),
.W_3(W_3_x427),
.W_4(W_4_x427),
.W_5(W_5_x427),
.W_6(W_6_x427),
.W_7(W_7_x427),
.W_8(W_8_x427),
.W_9(W_9_x427)
) u_28X28_x427 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x427),
 .score_0 (score_0_x427),
 .score_1 (score_1_x427),
 .score_2 (score_2_x427),
 .score_3 (score_3_x427),
 .score_4 (score_4_x427),
 .score_5 (score_5_x427),
 .score_6 (score_6_x427),
 .score_7 (score_7_x427),
 .score_8 (score_8_x427),
 .score_9 (score_9_x427)
);
 
myram_28X28 #(
.ID(428),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x428),
.W_1(W_1_x428),
.W_2(W_2_x428),
.W_3(W_3_x428),
.W_4(W_4_x428),
.W_5(W_5_x428),
.W_6(W_6_x428),
.W_7(W_7_x428),
.W_8(W_8_x428),
.W_9(W_9_x428)
) u_28X28_x428 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x428),
 .score_0 (score_0_x428),
 .score_1 (score_1_x428),
 .score_2 (score_2_x428),
 .score_3 (score_3_x428),
 .score_4 (score_4_x428),
 .score_5 (score_5_x428),
 .score_6 (score_6_x428),
 .score_7 (score_7_x428),
 .score_8 (score_8_x428),
 .score_9 (score_9_x428)
);
 
myram_28X28 #(
.ID(429),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x429),
.W_1(W_1_x429),
.W_2(W_2_x429),
.W_3(W_3_x429),
.W_4(W_4_x429),
.W_5(W_5_x429),
.W_6(W_6_x429),
.W_7(W_7_x429),
.W_8(W_8_x429),
.W_9(W_9_x429)
) u_28X28_x429 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x429),
 .score_0 (score_0_x429),
 .score_1 (score_1_x429),
 .score_2 (score_2_x429),
 .score_3 (score_3_x429),
 .score_4 (score_4_x429),
 .score_5 (score_5_x429),
 .score_6 (score_6_x429),
 .score_7 (score_7_x429),
 .score_8 (score_8_x429),
 .score_9 (score_9_x429)
);
 
myram_28X28 #(
.ID(430),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x430),
.W_1(W_1_x430),
.W_2(W_2_x430),
.W_3(W_3_x430),
.W_4(W_4_x430),
.W_5(W_5_x430),
.W_6(W_6_x430),
.W_7(W_7_x430),
.W_8(W_8_x430),
.W_9(W_9_x430)
) u_28X28_x430 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x430),
 .score_0 (score_0_x430),
 .score_1 (score_1_x430),
 .score_2 (score_2_x430),
 .score_3 (score_3_x430),
 .score_4 (score_4_x430),
 .score_5 (score_5_x430),
 .score_6 (score_6_x430),
 .score_7 (score_7_x430),
 .score_8 (score_8_x430),
 .score_9 (score_9_x430)
);
 
myram_28X28 #(
.ID(431),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x431),
.W_1(W_1_x431),
.W_2(W_2_x431),
.W_3(W_3_x431),
.W_4(W_4_x431),
.W_5(W_5_x431),
.W_6(W_6_x431),
.W_7(W_7_x431),
.W_8(W_8_x431),
.W_9(W_9_x431)
) u_28X28_x431 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x431),
 .score_0 (score_0_x431),
 .score_1 (score_1_x431),
 .score_2 (score_2_x431),
 .score_3 (score_3_x431),
 .score_4 (score_4_x431),
 .score_5 (score_5_x431),
 .score_6 (score_6_x431),
 .score_7 (score_7_x431),
 .score_8 (score_8_x431),
 .score_9 (score_9_x431)
);
 
myram_28X28 #(
.ID(432),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x432),
.W_1(W_1_x432),
.W_2(W_2_x432),
.W_3(W_3_x432),
.W_4(W_4_x432),
.W_5(W_5_x432),
.W_6(W_6_x432),
.W_7(W_7_x432),
.W_8(W_8_x432),
.W_9(W_9_x432)
) u_28X28_x432 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x432),
 .score_0 (score_0_x432),
 .score_1 (score_1_x432),
 .score_2 (score_2_x432),
 .score_3 (score_3_x432),
 .score_4 (score_4_x432),
 .score_5 (score_5_x432),
 .score_6 (score_6_x432),
 .score_7 (score_7_x432),
 .score_8 (score_8_x432),
 .score_9 (score_9_x432)
);
 
myram_28X28 #(
.ID(433),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x433),
.W_1(W_1_x433),
.W_2(W_2_x433),
.W_3(W_3_x433),
.W_4(W_4_x433),
.W_5(W_5_x433),
.W_6(W_6_x433),
.W_7(W_7_x433),
.W_8(W_8_x433),
.W_9(W_9_x433)
) u_28X28_x433 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x433),
 .score_0 (score_0_x433),
 .score_1 (score_1_x433),
 .score_2 (score_2_x433),
 .score_3 (score_3_x433),
 .score_4 (score_4_x433),
 .score_5 (score_5_x433),
 .score_6 (score_6_x433),
 .score_7 (score_7_x433),
 .score_8 (score_8_x433),
 .score_9 (score_9_x433)
);
 
myram_28X28 #(
.ID(434),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x434),
.W_1(W_1_x434),
.W_2(W_2_x434),
.W_3(W_3_x434),
.W_4(W_4_x434),
.W_5(W_5_x434),
.W_6(W_6_x434),
.W_7(W_7_x434),
.W_8(W_8_x434),
.W_9(W_9_x434)
) u_28X28_x434 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x434),
 .score_0 (score_0_x434),
 .score_1 (score_1_x434),
 .score_2 (score_2_x434),
 .score_3 (score_3_x434),
 .score_4 (score_4_x434),
 .score_5 (score_5_x434),
 .score_6 (score_6_x434),
 .score_7 (score_7_x434),
 .score_8 (score_8_x434),
 .score_9 (score_9_x434)
);
 
myram_28X28 #(
.ID(435),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x435),
.W_1(W_1_x435),
.W_2(W_2_x435),
.W_3(W_3_x435),
.W_4(W_4_x435),
.W_5(W_5_x435),
.W_6(W_6_x435),
.W_7(W_7_x435),
.W_8(W_8_x435),
.W_9(W_9_x435)
) u_28X28_x435 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x435),
 .score_0 (score_0_x435),
 .score_1 (score_1_x435),
 .score_2 (score_2_x435),
 .score_3 (score_3_x435),
 .score_4 (score_4_x435),
 .score_5 (score_5_x435),
 .score_6 (score_6_x435),
 .score_7 (score_7_x435),
 .score_8 (score_8_x435),
 .score_9 (score_9_x435)
);
 
myram_28X28 #(
.ID(436),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x436),
.W_1(W_1_x436),
.W_2(W_2_x436),
.W_3(W_3_x436),
.W_4(W_4_x436),
.W_5(W_5_x436),
.W_6(W_6_x436),
.W_7(W_7_x436),
.W_8(W_8_x436),
.W_9(W_9_x436)
) u_28X28_x436 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x436),
 .score_0 (score_0_x436),
 .score_1 (score_1_x436),
 .score_2 (score_2_x436),
 .score_3 (score_3_x436),
 .score_4 (score_4_x436),
 .score_5 (score_5_x436),
 .score_6 (score_6_x436),
 .score_7 (score_7_x436),
 .score_8 (score_8_x436),
 .score_9 (score_9_x436)
);
 
myram_28X28 #(
.ID(437),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x437),
.W_1(W_1_x437),
.W_2(W_2_x437),
.W_3(W_3_x437),
.W_4(W_4_x437),
.W_5(W_5_x437),
.W_6(W_6_x437),
.W_7(W_7_x437),
.W_8(W_8_x437),
.W_9(W_9_x437)
) u_28X28_x437 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x437),
 .score_0 (score_0_x437),
 .score_1 (score_1_x437),
 .score_2 (score_2_x437),
 .score_3 (score_3_x437),
 .score_4 (score_4_x437),
 .score_5 (score_5_x437),
 .score_6 (score_6_x437),
 .score_7 (score_7_x437),
 .score_8 (score_8_x437),
 .score_9 (score_9_x437)
);
 
myram_28X28 #(
.ID(438),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x438),
.W_1(W_1_x438),
.W_2(W_2_x438),
.W_3(W_3_x438),
.W_4(W_4_x438),
.W_5(W_5_x438),
.W_6(W_6_x438),
.W_7(W_7_x438),
.W_8(W_8_x438),
.W_9(W_9_x438)
) u_28X28_x438 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x438),
 .score_0 (score_0_x438),
 .score_1 (score_1_x438),
 .score_2 (score_2_x438),
 .score_3 (score_3_x438),
 .score_4 (score_4_x438),
 .score_5 (score_5_x438),
 .score_6 (score_6_x438),
 .score_7 (score_7_x438),
 .score_8 (score_8_x438),
 .score_9 (score_9_x438)
);
 
myram_28X28 #(
.ID(439),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x439),
.W_1(W_1_x439),
.W_2(W_2_x439),
.W_3(W_3_x439),
.W_4(W_4_x439),
.W_5(W_5_x439),
.W_6(W_6_x439),
.W_7(W_7_x439),
.W_8(W_8_x439),
.W_9(W_9_x439)
) u_28X28_x439 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x439),
 .score_0 (score_0_x439),
 .score_1 (score_1_x439),
 .score_2 (score_2_x439),
 .score_3 (score_3_x439),
 .score_4 (score_4_x439),
 .score_5 (score_5_x439),
 .score_6 (score_6_x439),
 .score_7 (score_7_x439),
 .score_8 (score_8_x439),
 .score_9 (score_9_x439)
);
 
myram_28X28 #(
.ID(440),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x440),
.W_1(W_1_x440),
.W_2(W_2_x440),
.W_3(W_3_x440),
.W_4(W_4_x440),
.W_5(W_5_x440),
.W_6(W_6_x440),
.W_7(W_7_x440),
.W_8(W_8_x440),
.W_9(W_9_x440)
) u_28X28_x440 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x440),
 .score_0 (score_0_x440),
 .score_1 (score_1_x440),
 .score_2 (score_2_x440),
 .score_3 (score_3_x440),
 .score_4 (score_4_x440),
 .score_5 (score_5_x440),
 .score_6 (score_6_x440),
 .score_7 (score_7_x440),
 .score_8 (score_8_x440),
 .score_9 (score_9_x440)
);
 
myram_28X28 #(
.ID(441),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x441),
.W_1(W_1_x441),
.W_2(W_2_x441),
.W_3(W_3_x441),
.W_4(W_4_x441),
.W_5(W_5_x441),
.W_6(W_6_x441),
.W_7(W_7_x441),
.W_8(W_8_x441),
.W_9(W_9_x441)
) u_28X28_x441 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x441),
 .score_0 (score_0_x441),
 .score_1 (score_1_x441),
 .score_2 (score_2_x441),
 .score_3 (score_3_x441),
 .score_4 (score_4_x441),
 .score_5 (score_5_x441),
 .score_6 (score_6_x441),
 .score_7 (score_7_x441),
 .score_8 (score_8_x441),
 .score_9 (score_9_x441)
);
 
myram_28X28 #(
.ID(442),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x442),
.W_1(W_1_x442),
.W_2(W_2_x442),
.W_3(W_3_x442),
.W_4(W_4_x442),
.W_5(W_5_x442),
.W_6(W_6_x442),
.W_7(W_7_x442),
.W_8(W_8_x442),
.W_9(W_9_x442)
) u_28X28_x442 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x442),
 .score_0 (score_0_x442),
 .score_1 (score_1_x442),
 .score_2 (score_2_x442),
 .score_3 (score_3_x442),
 .score_4 (score_4_x442),
 .score_5 (score_5_x442),
 .score_6 (score_6_x442),
 .score_7 (score_7_x442),
 .score_8 (score_8_x442),
 .score_9 (score_9_x442)
);
 
myram_28X28 #(
.ID(443),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x443),
.W_1(W_1_x443),
.W_2(W_2_x443),
.W_3(W_3_x443),
.W_4(W_4_x443),
.W_5(W_5_x443),
.W_6(W_6_x443),
.W_7(W_7_x443),
.W_8(W_8_x443),
.W_9(W_9_x443)
) u_28X28_x443 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x443),
 .score_0 (score_0_x443),
 .score_1 (score_1_x443),
 .score_2 (score_2_x443),
 .score_3 (score_3_x443),
 .score_4 (score_4_x443),
 .score_5 (score_5_x443),
 .score_6 (score_6_x443),
 .score_7 (score_7_x443),
 .score_8 (score_8_x443),
 .score_9 (score_9_x443)
);
 
myram_28X28 #(
.ID(444),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x444),
.W_1(W_1_x444),
.W_2(W_2_x444),
.W_3(W_3_x444),
.W_4(W_4_x444),
.W_5(W_5_x444),
.W_6(W_6_x444),
.W_7(W_7_x444),
.W_8(W_8_x444),
.W_9(W_9_x444)
) u_28X28_x444 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x444),
 .score_0 (score_0_x444),
 .score_1 (score_1_x444),
 .score_2 (score_2_x444),
 .score_3 (score_3_x444),
 .score_4 (score_4_x444),
 .score_5 (score_5_x444),
 .score_6 (score_6_x444),
 .score_7 (score_7_x444),
 .score_8 (score_8_x444),
 .score_9 (score_9_x444)
);
 
myram_28X28 #(
.ID(445),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x445),
.W_1(W_1_x445),
.W_2(W_2_x445),
.W_3(W_3_x445),
.W_4(W_4_x445),
.W_5(W_5_x445),
.W_6(W_6_x445),
.W_7(W_7_x445),
.W_8(W_8_x445),
.W_9(W_9_x445)
) u_28X28_x445 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x445),
 .score_0 (score_0_x445),
 .score_1 (score_1_x445),
 .score_2 (score_2_x445),
 .score_3 (score_3_x445),
 .score_4 (score_4_x445),
 .score_5 (score_5_x445),
 .score_6 (score_6_x445),
 .score_7 (score_7_x445),
 .score_8 (score_8_x445),
 .score_9 (score_9_x445)
);
 
myram_28X28 #(
.ID(446),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x446),
.W_1(W_1_x446),
.W_2(W_2_x446),
.W_3(W_3_x446),
.W_4(W_4_x446),
.W_5(W_5_x446),
.W_6(W_6_x446),
.W_7(W_7_x446),
.W_8(W_8_x446),
.W_9(W_9_x446)
) u_28X28_x446 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x446),
 .score_0 (score_0_x446),
 .score_1 (score_1_x446),
 .score_2 (score_2_x446),
 .score_3 (score_3_x446),
 .score_4 (score_4_x446),
 .score_5 (score_5_x446),
 .score_6 (score_6_x446),
 .score_7 (score_7_x446),
 .score_8 (score_8_x446),
 .score_9 (score_9_x446)
);
 
myram_28X28 #(
.ID(447),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x447),
.W_1(W_1_x447),
.W_2(W_2_x447),
.W_3(W_3_x447),
.W_4(W_4_x447),
.W_5(W_5_x447),
.W_6(W_6_x447),
.W_7(W_7_x447),
.W_8(W_8_x447),
.W_9(W_9_x447)
) u_28X28_x447 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x447),
 .score_0 (score_0_x447),
 .score_1 (score_1_x447),
 .score_2 (score_2_x447),
 .score_3 (score_3_x447),
 .score_4 (score_4_x447),
 .score_5 (score_5_x447),
 .score_6 (score_6_x447),
 .score_7 (score_7_x447),
 .score_8 (score_8_x447),
 .score_9 (score_9_x447)
);
 
myram_28X28 #(
.ID(448),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x448),
.W_1(W_1_x448),
.W_2(W_2_x448),
.W_3(W_3_x448),
.W_4(W_4_x448),
.W_5(W_5_x448),
.W_6(W_6_x448),
.W_7(W_7_x448),
.W_8(W_8_x448),
.W_9(W_9_x448)
) u_28X28_x448 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x448),
 .score_0 (score_0_x448),
 .score_1 (score_1_x448),
 .score_2 (score_2_x448),
 .score_3 (score_3_x448),
 .score_4 (score_4_x448),
 .score_5 (score_5_x448),
 .score_6 (score_6_x448),
 .score_7 (score_7_x448),
 .score_8 (score_8_x448),
 .score_9 (score_9_x448)
);
 
myram_28X28 #(
.ID(449),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x449),
.W_1(W_1_x449),
.W_2(W_2_x449),
.W_3(W_3_x449),
.W_4(W_4_x449),
.W_5(W_5_x449),
.W_6(W_6_x449),
.W_7(W_7_x449),
.W_8(W_8_x449),
.W_9(W_9_x449)
) u_28X28_x449 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x449),
 .score_0 (score_0_x449),
 .score_1 (score_1_x449),
 .score_2 (score_2_x449),
 .score_3 (score_3_x449),
 .score_4 (score_4_x449),
 .score_5 (score_5_x449),
 .score_6 (score_6_x449),
 .score_7 (score_7_x449),
 .score_8 (score_8_x449),
 .score_9 (score_9_x449)
);
 
myram_28X28 #(
.ID(450),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x450),
.W_1(W_1_x450),
.W_2(W_2_x450),
.W_3(W_3_x450),
.W_4(W_4_x450),
.W_5(W_5_x450),
.W_6(W_6_x450),
.W_7(W_7_x450),
.W_8(W_8_x450),
.W_9(W_9_x450)
) u_28X28_x450 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x450),
 .score_0 (score_0_x450),
 .score_1 (score_1_x450),
 .score_2 (score_2_x450),
 .score_3 (score_3_x450),
 .score_4 (score_4_x450),
 .score_5 (score_5_x450),
 .score_6 (score_6_x450),
 .score_7 (score_7_x450),
 .score_8 (score_8_x450),
 .score_9 (score_9_x450)
);
 
myram_28X28 #(
.ID(451),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x451),
.W_1(W_1_x451),
.W_2(W_2_x451),
.W_3(W_3_x451),
.W_4(W_4_x451),
.W_5(W_5_x451),
.W_6(W_6_x451),
.W_7(W_7_x451),
.W_8(W_8_x451),
.W_9(W_9_x451)
) u_28X28_x451 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x451),
 .score_0 (score_0_x451),
 .score_1 (score_1_x451),
 .score_2 (score_2_x451),
 .score_3 (score_3_x451),
 .score_4 (score_4_x451),
 .score_5 (score_5_x451),
 .score_6 (score_6_x451),
 .score_7 (score_7_x451),
 .score_8 (score_8_x451),
 .score_9 (score_9_x451)
);
 
myram_28X28 #(
.ID(452),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x452),
.W_1(W_1_x452),
.W_2(W_2_x452),
.W_3(W_3_x452),
.W_4(W_4_x452),
.W_5(W_5_x452),
.W_6(W_6_x452),
.W_7(W_7_x452),
.W_8(W_8_x452),
.W_9(W_9_x452)
) u_28X28_x452 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x452),
 .score_0 (score_0_x452),
 .score_1 (score_1_x452),
 .score_2 (score_2_x452),
 .score_3 (score_3_x452),
 .score_4 (score_4_x452),
 .score_5 (score_5_x452),
 .score_6 (score_6_x452),
 .score_7 (score_7_x452),
 .score_8 (score_8_x452),
 .score_9 (score_9_x452)
);
 
myram_28X28 #(
.ID(453),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x453),
.W_1(W_1_x453),
.W_2(W_2_x453),
.W_3(W_3_x453),
.W_4(W_4_x453),
.W_5(W_5_x453),
.W_6(W_6_x453),
.W_7(W_7_x453),
.W_8(W_8_x453),
.W_9(W_9_x453)
) u_28X28_x453 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x453),
 .score_0 (score_0_x453),
 .score_1 (score_1_x453),
 .score_2 (score_2_x453),
 .score_3 (score_3_x453),
 .score_4 (score_4_x453),
 .score_5 (score_5_x453),
 .score_6 (score_6_x453),
 .score_7 (score_7_x453),
 .score_8 (score_8_x453),
 .score_9 (score_9_x453)
);
 
myram_28X28 #(
.ID(454),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x454),
.W_1(W_1_x454),
.W_2(W_2_x454),
.W_3(W_3_x454),
.W_4(W_4_x454),
.W_5(W_5_x454),
.W_6(W_6_x454),
.W_7(W_7_x454),
.W_8(W_8_x454),
.W_9(W_9_x454)
) u_28X28_x454 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x454),
 .score_0 (score_0_x454),
 .score_1 (score_1_x454),
 .score_2 (score_2_x454),
 .score_3 (score_3_x454),
 .score_4 (score_4_x454),
 .score_5 (score_5_x454),
 .score_6 (score_6_x454),
 .score_7 (score_7_x454),
 .score_8 (score_8_x454),
 .score_9 (score_9_x454)
);
 
myram_28X28 #(
.ID(455),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x455),
.W_1(W_1_x455),
.W_2(W_2_x455),
.W_3(W_3_x455),
.W_4(W_4_x455),
.W_5(W_5_x455),
.W_6(W_6_x455),
.W_7(W_7_x455),
.W_8(W_8_x455),
.W_9(W_9_x455)
) u_28X28_x455 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x455),
 .score_0 (score_0_x455),
 .score_1 (score_1_x455),
 .score_2 (score_2_x455),
 .score_3 (score_3_x455),
 .score_4 (score_4_x455),
 .score_5 (score_5_x455),
 .score_6 (score_6_x455),
 .score_7 (score_7_x455),
 .score_8 (score_8_x455),
 .score_9 (score_9_x455)
);
 
myram_28X28 #(
.ID(456),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x456),
.W_1(W_1_x456),
.W_2(W_2_x456),
.W_3(W_3_x456),
.W_4(W_4_x456),
.W_5(W_5_x456),
.W_6(W_6_x456),
.W_7(W_7_x456),
.W_8(W_8_x456),
.W_9(W_9_x456)
) u_28X28_x456 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x456),
 .score_0 (score_0_x456),
 .score_1 (score_1_x456),
 .score_2 (score_2_x456),
 .score_3 (score_3_x456),
 .score_4 (score_4_x456),
 .score_5 (score_5_x456),
 .score_6 (score_6_x456),
 .score_7 (score_7_x456),
 .score_8 (score_8_x456),
 .score_9 (score_9_x456)
);
 
myram_28X28 #(
.ID(457),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x457),
.W_1(W_1_x457),
.W_2(W_2_x457),
.W_3(W_3_x457),
.W_4(W_4_x457),
.W_5(W_5_x457),
.W_6(W_6_x457),
.W_7(W_7_x457),
.W_8(W_8_x457),
.W_9(W_9_x457)
) u_28X28_x457 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x457),
 .score_0 (score_0_x457),
 .score_1 (score_1_x457),
 .score_2 (score_2_x457),
 .score_3 (score_3_x457),
 .score_4 (score_4_x457),
 .score_5 (score_5_x457),
 .score_6 (score_6_x457),
 .score_7 (score_7_x457),
 .score_8 (score_8_x457),
 .score_9 (score_9_x457)
);
 
myram_28X28 #(
.ID(458),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x458),
.W_1(W_1_x458),
.W_2(W_2_x458),
.W_3(W_3_x458),
.W_4(W_4_x458),
.W_5(W_5_x458),
.W_6(W_6_x458),
.W_7(W_7_x458),
.W_8(W_8_x458),
.W_9(W_9_x458)
) u_28X28_x458 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x458),
 .score_0 (score_0_x458),
 .score_1 (score_1_x458),
 .score_2 (score_2_x458),
 .score_3 (score_3_x458),
 .score_4 (score_4_x458),
 .score_5 (score_5_x458),
 .score_6 (score_6_x458),
 .score_7 (score_7_x458),
 .score_8 (score_8_x458),
 .score_9 (score_9_x458)
);
 
myram_28X28 #(
.ID(459),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x459),
.W_1(W_1_x459),
.W_2(W_2_x459),
.W_3(W_3_x459),
.W_4(W_4_x459),
.W_5(W_5_x459),
.W_6(W_6_x459),
.W_7(W_7_x459),
.W_8(W_8_x459),
.W_9(W_9_x459)
) u_28X28_x459 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x459),
 .score_0 (score_0_x459),
 .score_1 (score_1_x459),
 .score_2 (score_2_x459),
 .score_3 (score_3_x459),
 .score_4 (score_4_x459),
 .score_5 (score_5_x459),
 .score_6 (score_6_x459),
 .score_7 (score_7_x459),
 .score_8 (score_8_x459),
 .score_9 (score_9_x459)
);
 
myram_28X28 #(
.ID(460),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x460),
.W_1(W_1_x460),
.W_2(W_2_x460),
.W_3(W_3_x460),
.W_4(W_4_x460),
.W_5(W_5_x460),
.W_6(W_6_x460),
.W_7(W_7_x460),
.W_8(W_8_x460),
.W_9(W_9_x460)
) u_28X28_x460 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x460),
 .score_0 (score_0_x460),
 .score_1 (score_1_x460),
 .score_2 (score_2_x460),
 .score_3 (score_3_x460),
 .score_4 (score_4_x460),
 .score_5 (score_5_x460),
 .score_6 (score_6_x460),
 .score_7 (score_7_x460),
 .score_8 (score_8_x460),
 .score_9 (score_9_x460)
);
 
myram_28X28 #(
.ID(461),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x461),
.W_1(W_1_x461),
.W_2(W_2_x461),
.W_3(W_3_x461),
.W_4(W_4_x461),
.W_5(W_5_x461),
.W_6(W_6_x461),
.W_7(W_7_x461),
.W_8(W_8_x461),
.W_9(W_9_x461)
) u_28X28_x461 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x461),
 .score_0 (score_0_x461),
 .score_1 (score_1_x461),
 .score_2 (score_2_x461),
 .score_3 (score_3_x461),
 .score_4 (score_4_x461),
 .score_5 (score_5_x461),
 .score_6 (score_6_x461),
 .score_7 (score_7_x461),
 .score_8 (score_8_x461),
 .score_9 (score_9_x461)
);
 
myram_28X28 #(
.ID(462),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x462),
.W_1(W_1_x462),
.W_2(W_2_x462),
.W_3(W_3_x462),
.W_4(W_4_x462),
.W_5(W_5_x462),
.W_6(W_6_x462),
.W_7(W_7_x462),
.W_8(W_8_x462),
.W_9(W_9_x462)
) u_28X28_x462 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x462),
 .score_0 (score_0_x462),
 .score_1 (score_1_x462),
 .score_2 (score_2_x462),
 .score_3 (score_3_x462),
 .score_4 (score_4_x462),
 .score_5 (score_5_x462),
 .score_6 (score_6_x462),
 .score_7 (score_7_x462),
 .score_8 (score_8_x462),
 .score_9 (score_9_x462)
);
 
myram_28X28 #(
.ID(463),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x463),
.W_1(W_1_x463),
.W_2(W_2_x463),
.W_3(W_3_x463),
.W_4(W_4_x463),
.W_5(W_5_x463),
.W_6(W_6_x463),
.W_7(W_7_x463),
.W_8(W_8_x463),
.W_9(W_9_x463)
) u_28X28_x463 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x463),
 .score_0 (score_0_x463),
 .score_1 (score_1_x463),
 .score_2 (score_2_x463),
 .score_3 (score_3_x463),
 .score_4 (score_4_x463),
 .score_5 (score_5_x463),
 .score_6 (score_6_x463),
 .score_7 (score_7_x463),
 .score_8 (score_8_x463),
 .score_9 (score_9_x463)
);
 
myram_28X28 #(
.ID(464),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x464),
.W_1(W_1_x464),
.W_2(W_2_x464),
.W_3(W_3_x464),
.W_4(W_4_x464),
.W_5(W_5_x464),
.W_6(W_6_x464),
.W_7(W_7_x464),
.W_8(W_8_x464),
.W_9(W_9_x464)
) u_28X28_x464 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x464),
 .score_0 (score_0_x464),
 .score_1 (score_1_x464),
 .score_2 (score_2_x464),
 .score_3 (score_3_x464),
 .score_4 (score_4_x464),
 .score_5 (score_5_x464),
 .score_6 (score_6_x464),
 .score_7 (score_7_x464),
 .score_8 (score_8_x464),
 .score_9 (score_9_x464)
);
 
myram_28X28 #(
.ID(465),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x465),
.W_1(W_1_x465),
.W_2(W_2_x465),
.W_3(W_3_x465),
.W_4(W_4_x465),
.W_5(W_5_x465),
.W_6(W_6_x465),
.W_7(W_7_x465),
.W_8(W_8_x465),
.W_9(W_9_x465)
) u_28X28_x465 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x465),
 .score_0 (score_0_x465),
 .score_1 (score_1_x465),
 .score_2 (score_2_x465),
 .score_3 (score_3_x465),
 .score_4 (score_4_x465),
 .score_5 (score_5_x465),
 .score_6 (score_6_x465),
 .score_7 (score_7_x465),
 .score_8 (score_8_x465),
 .score_9 (score_9_x465)
);
 
myram_28X28 #(
.ID(466),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x466),
.W_1(W_1_x466),
.W_2(W_2_x466),
.W_3(W_3_x466),
.W_4(W_4_x466),
.W_5(W_5_x466),
.W_6(W_6_x466),
.W_7(W_7_x466),
.W_8(W_8_x466),
.W_9(W_9_x466)
) u_28X28_x466 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x466),
 .score_0 (score_0_x466),
 .score_1 (score_1_x466),
 .score_2 (score_2_x466),
 .score_3 (score_3_x466),
 .score_4 (score_4_x466),
 .score_5 (score_5_x466),
 .score_6 (score_6_x466),
 .score_7 (score_7_x466),
 .score_8 (score_8_x466),
 .score_9 (score_9_x466)
);
 
myram_28X28 #(
.ID(467),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x467),
.W_1(W_1_x467),
.W_2(W_2_x467),
.W_3(W_3_x467),
.W_4(W_4_x467),
.W_5(W_5_x467),
.W_6(W_6_x467),
.W_7(W_7_x467),
.W_8(W_8_x467),
.W_9(W_9_x467)
) u_28X28_x467 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x467),
 .score_0 (score_0_x467),
 .score_1 (score_1_x467),
 .score_2 (score_2_x467),
 .score_3 (score_3_x467),
 .score_4 (score_4_x467),
 .score_5 (score_5_x467),
 .score_6 (score_6_x467),
 .score_7 (score_7_x467),
 .score_8 (score_8_x467),
 .score_9 (score_9_x467)
);
 
myram_28X28 #(
.ID(468),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x468),
.W_1(W_1_x468),
.W_2(W_2_x468),
.W_3(W_3_x468),
.W_4(W_4_x468),
.W_5(W_5_x468),
.W_6(W_6_x468),
.W_7(W_7_x468),
.W_8(W_8_x468),
.W_9(W_9_x468)
) u_28X28_x468 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x468),
 .score_0 (score_0_x468),
 .score_1 (score_1_x468),
 .score_2 (score_2_x468),
 .score_3 (score_3_x468),
 .score_4 (score_4_x468),
 .score_5 (score_5_x468),
 .score_6 (score_6_x468),
 .score_7 (score_7_x468),
 .score_8 (score_8_x468),
 .score_9 (score_9_x468)
);
 
myram_28X28 #(
.ID(469),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x469),
.W_1(W_1_x469),
.W_2(W_2_x469),
.W_3(W_3_x469),
.W_4(W_4_x469),
.W_5(W_5_x469),
.W_6(W_6_x469),
.W_7(W_7_x469),
.W_8(W_8_x469),
.W_9(W_9_x469)
) u_28X28_x469 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x469),
 .score_0 (score_0_x469),
 .score_1 (score_1_x469),
 .score_2 (score_2_x469),
 .score_3 (score_3_x469),
 .score_4 (score_4_x469),
 .score_5 (score_5_x469),
 .score_6 (score_6_x469),
 .score_7 (score_7_x469),
 .score_8 (score_8_x469),
 .score_9 (score_9_x469)
);
 
myram_28X28 #(
.ID(470),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x470),
.W_1(W_1_x470),
.W_2(W_2_x470),
.W_3(W_3_x470),
.W_4(W_4_x470),
.W_5(W_5_x470),
.W_6(W_6_x470),
.W_7(W_7_x470),
.W_8(W_8_x470),
.W_9(W_9_x470)
) u_28X28_x470 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x470),
 .score_0 (score_0_x470),
 .score_1 (score_1_x470),
 .score_2 (score_2_x470),
 .score_3 (score_3_x470),
 .score_4 (score_4_x470),
 .score_5 (score_5_x470),
 .score_6 (score_6_x470),
 .score_7 (score_7_x470),
 .score_8 (score_8_x470),
 .score_9 (score_9_x470)
);
 
myram_28X28 #(
.ID(471),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x471),
.W_1(W_1_x471),
.W_2(W_2_x471),
.W_3(W_3_x471),
.W_4(W_4_x471),
.W_5(W_5_x471),
.W_6(W_6_x471),
.W_7(W_7_x471),
.W_8(W_8_x471),
.W_9(W_9_x471)
) u_28X28_x471 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x471),
 .score_0 (score_0_x471),
 .score_1 (score_1_x471),
 .score_2 (score_2_x471),
 .score_3 (score_3_x471),
 .score_4 (score_4_x471),
 .score_5 (score_5_x471),
 .score_6 (score_6_x471),
 .score_7 (score_7_x471),
 .score_8 (score_8_x471),
 .score_9 (score_9_x471)
);
 
myram_28X28 #(
.ID(472),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x472),
.W_1(W_1_x472),
.W_2(W_2_x472),
.W_3(W_3_x472),
.W_4(W_4_x472),
.W_5(W_5_x472),
.W_6(W_6_x472),
.W_7(W_7_x472),
.W_8(W_8_x472),
.W_9(W_9_x472)
) u_28X28_x472 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x472),
 .score_0 (score_0_x472),
 .score_1 (score_1_x472),
 .score_2 (score_2_x472),
 .score_3 (score_3_x472),
 .score_4 (score_4_x472),
 .score_5 (score_5_x472),
 .score_6 (score_6_x472),
 .score_7 (score_7_x472),
 .score_8 (score_8_x472),
 .score_9 (score_9_x472)
);
 
myram_28X28 #(
.ID(473),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x473),
.W_1(W_1_x473),
.W_2(W_2_x473),
.W_3(W_3_x473),
.W_4(W_4_x473),
.W_5(W_5_x473),
.W_6(W_6_x473),
.W_7(W_7_x473),
.W_8(W_8_x473),
.W_9(W_9_x473)
) u_28X28_x473 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x473),
 .score_0 (score_0_x473),
 .score_1 (score_1_x473),
 .score_2 (score_2_x473),
 .score_3 (score_3_x473),
 .score_4 (score_4_x473),
 .score_5 (score_5_x473),
 .score_6 (score_6_x473),
 .score_7 (score_7_x473),
 .score_8 (score_8_x473),
 .score_9 (score_9_x473)
);
 
myram_28X28 #(
.ID(474),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x474),
.W_1(W_1_x474),
.W_2(W_2_x474),
.W_3(W_3_x474),
.W_4(W_4_x474),
.W_5(W_5_x474),
.W_6(W_6_x474),
.W_7(W_7_x474),
.W_8(W_8_x474),
.W_9(W_9_x474)
) u_28X28_x474 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x474),
 .score_0 (score_0_x474),
 .score_1 (score_1_x474),
 .score_2 (score_2_x474),
 .score_3 (score_3_x474),
 .score_4 (score_4_x474),
 .score_5 (score_5_x474),
 .score_6 (score_6_x474),
 .score_7 (score_7_x474),
 .score_8 (score_8_x474),
 .score_9 (score_9_x474)
);
 
myram_28X28 #(
.ID(475),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x475),
.W_1(W_1_x475),
.W_2(W_2_x475),
.W_3(W_3_x475),
.W_4(W_4_x475),
.W_5(W_5_x475),
.W_6(W_6_x475),
.W_7(W_7_x475),
.W_8(W_8_x475),
.W_9(W_9_x475)
) u_28X28_x475 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x475),
 .score_0 (score_0_x475),
 .score_1 (score_1_x475),
 .score_2 (score_2_x475),
 .score_3 (score_3_x475),
 .score_4 (score_4_x475),
 .score_5 (score_5_x475),
 .score_6 (score_6_x475),
 .score_7 (score_7_x475),
 .score_8 (score_8_x475),
 .score_9 (score_9_x475)
);
 
myram_28X28 #(
.ID(476),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x476),
.W_1(W_1_x476),
.W_2(W_2_x476),
.W_3(W_3_x476),
.W_4(W_4_x476),
.W_5(W_5_x476),
.W_6(W_6_x476),
.W_7(W_7_x476),
.W_8(W_8_x476),
.W_9(W_9_x476)
) u_28X28_x476 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x476),
 .score_0 (score_0_x476),
 .score_1 (score_1_x476),
 .score_2 (score_2_x476),
 .score_3 (score_3_x476),
 .score_4 (score_4_x476),
 .score_5 (score_5_x476),
 .score_6 (score_6_x476),
 .score_7 (score_7_x476),
 .score_8 (score_8_x476),
 .score_9 (score_9_x476)
);
 
myram_28X28 #(
.ID(477),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x477),
.W_1(W_1_x477),
.W_2(W_2_x477),
.W_3(W_3_x477),
.W_4(W_4_x477),
.W_5(W_5_x477),
.W_6(W_6_x477),
.W_7(W_7_x477),
.W_8(W_8_x477),
.W_9(W_9_x477)
) u_28X28_x477 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x477),
 .score_0 (score_0_x477),
 .score_1 (score_1_x477),
 .score_2 (score_2_x477),
 .score_3 (score_3_x477),
 .score_4 (score_4_x477),
 .score_5 (score_5_x477),
 .score_6 (score_6_x477),
 .score_7 (score_7_x477),
 .score_8 (score_8_x477),
 .score_9 (score_9_x477)
);
 
myram_28X28 #(
.ID(478),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x478),
.W_1(W_1_x478),
.W_2(W_2_x478),
.W_3(W_3_x478),
.W_4(W_4_x478),
.W_5(W_5_x478),
.W_6(W_6_x478),
.W_7(W_7_x478),
.W_8(W_8_x478),
.W_9(W_9_x478)
) u_28X28_x478 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x478),
 .score_0 (score_0_x478),
 .score_1 (score_1_x478),
 .score_2 (score_2_x478),
 .score_3 (score_3_x478),
 .score_4 (score_4_x478),
 .score_5 (score_5_x478),
 .score_6 (score_6_x478),
 .score_7 (score_7_x478),
 .score_8 (score_8_x478),
 .score_9 (score_9_x478)
);
 
myram_28X28 #(
.ID(479),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x479),
.W_1(W_1_x479),
.W_2(W_2_x479),
.W_3(W_3_x479),
.W_4(W_4_x479),
.W_5(W_5_x479),
.W_6(W_6_x479),
.W_7(W_7_x479),
.W_8(W_8_x479),
.W_9(W_9_x479)
) u_28X28_x479 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x479),
 .score_0 (score_0_x479),
 .score_1 (score_1_x479),
 .score_2 (score_2_x479),
 .score_3 (score_3_x479),
 .score_4 (score_4_x479),
 .score_5 (score_5_x479),
 .score_6 (score_6_x479),
 .score_7 (score_7_x479),
 .score_8 (score_8_x479),
 .score_9 (score_9_x479)
);
 
myram_28X28 #(
.ID(480),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x480),
.W_1(W_1_x480),
.W_2(W_2_x480),
.W_3(W_3_x480),
.W_4(W_4_x480),
.W_5(W_5_x480),
.W_6(W_6_x480),
.W_7(W_7_x480),
.W_8(W_8_x480),
.W_9(W_9_x480)
) u_28X28_x480 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x480),
 .score_0 (score_0_x480),
 .score_1 (score_1_x480),
 .score_2 (score_2_x480),
 .score_3 (score_3_x480),
 .score_4 (score_4_x480),
 .score_5 (score_5_x480),
 .score_6 (score_6_x480),
 .score_7 (score_7_x480),
 .score_8 (score_8_x480),
 .score_9 (score_9_x480)
);
 
myram_28X28 #(
.ID(481),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x481),
.W_1(W_1_x481),
.W_2(W_2_x481),
.W_3(W_3_x481),
.W_4(W_4_x481),
.W_5(W_5_x481),
.W_6(W_6_x481),
.W_7(W_7_x481),
.W_8(W_8_x481),
.W_9(W_9_x481)
) u_28X28_x481 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x481),
 .score_0 (score_0_x481),
 .score_1 (score_1_x481),
 .score_2 (score_2_x481),
 .score_3 (score_3_x481),
 .score_4 (score_4_x481),
 .score_5 (score_5_x481),
 .score_6 (score_6_x481),
 .score_7 (score_7_x481),
 .score_8 (score_8_x481),
 .score_9 (score_9_x481)
);
 
myram_28X28 #(
.ID(482),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x482),
.W_1(W_1_x482),
.W_2(W_2_x482),
.W_3(W_3_x482),
.W_4(W_4_x482),
.W_5(W_5_x482),
.W_6(W_6_x482),
.W_7(W_7_x482),
.W_8(W_8_x482),
.W_9(W_9_x482)
) u_28X28_x482 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x482),
 .score_0 (score_0_x482),
 .score_1 (score_1_x482),
 .score_2 (score_2_x482),
 .score_3 (score_3_x482),
 .score_4 (score_4_x482),
 .score_5 (score_5_x482),
 .score_6 (score_6_x482),
 .score_7 (score_7_x482),
 .score_8 (score_8_x482),
 .score_9 (score_9_x482)
);
 
myram_28X28 #(
.ID(483),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x483),
.W_1(W_1_x483),
.W_2(W_2_x483),
.W_3(W_3_x483),
.W_4(W_4_x483),
.W_5(W_5_x483),
.W_6(W_6_x483),
.W_7(W_7_x483),
.W_8(W_8_x483),
.W_9(W_9_x483)
) u_28X28_x483 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x483),
 .score_0 (score_0_x483),
 .score_1 (score_1_x483),
 .score_2 (score_2_x483),
 .score_3 (score_3_x483),
 .score_4 (score_4_x483),
 .score_5 (score_5_x483),
 .score_6 (score_6_x483),
 .score_7 (score_7_x483),
 .score_8 (score_8_x483),
 .score_9 (score_9_x483)
);
 
myram_28X28 #(
.ID(484),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x484),
.W_1(W_1_x484),
.W_2(W_2_x484),
.W_3(W_3_x484),
.W_4(W_4_x484),
.W_5(W_5_x484),
.W_6(W_6_x484),
.W_7(W_7_x484),
.W_8(W_8_x484),
.W_9(W_9_x484)
) u_28X28_x484 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x484),
 .score_0 (score_0_x484),
 .score_1 (score_1_x484),
 .score_2 (score_2_x484),
 .score_3 (score_3_x484),
 .score_4 (score_4_x484),
 .score_5 (score_5_x484),
 .score_6 (score_6_x484),
 .score_7 (score_7_x484),
 .score_8 (score_8_x484),
 .score_9 (score_9_x484)
);
 
myram_28X28 #(
.ID(485),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x485),
.W_1(W_1_x485),
.W_2(W_2_x485),
.W_3(W_3_x485),
.W_4(W_4_x485),
.W_5(W_5_x485),
.W_6(W_6_x485),
.W_7(W_7_x485),
.W_8(W_8_x485),
.W_9(W_9_x485)
) u_28X28_x485 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x485),
 .score_0 (score_0_x485),
 .score_1 (score_1_x485),
 .score_2 (score_2_x485),
 .score_3 (score_3_x485),
 .score_4 (score_4_x485),
 .score_5 (score_5_x485),
 .score_6 (score_6_x485),
 .score_7 (score_7_x485),
 .score_8 (score_8_x485),
 .score_9 (score_9_x485)
);
 
myram_28X28 #(
.ID(486),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x486),
.W_1(W_1_x486),
.W_2(W_2_x486),
.W_3(W_3_x486),
.W_4(W_4_x486),
.W_5(W_5_x486),
.W_6(W_6_x486),
.W_7(W_7_x486),
.W_8(W_8_x486),
.W_9(W_9_x486)
) u_28X28_x486 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x486),
 .score_0 (score_0_x486),
 .score_1 (score_1_x486),
 .score_2 (score_2_x486),
 .score_3 (score_3_x486),
 .score_4 (score_4_x486),
 .score_5 (score_5_x486),
 .score_6 (score_6_x486),
 .score_7 (score_7_x486),
 .score_8 (score_8_x486),
 .score_9 (score_9_x486)
);
 
myram_28X28 #(
.ID(487),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x487),
.W_1(W_1_x487),
.W_2(W_2_x487),
.W_3(W_3_x487),
.W_4(W_4_x487),
.W_5(W_5_x487),
.W_6(W_6_x487),
.W_7(W_7_x487),
.W_8(W_8_x487),
.W_9(W_9_x487)
) u_28X28_x487 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x487),
 .score_0 (score_0_x487),
 .score_1 (score_1_x487),
 .score_2 (score_2_x487),
 .score_3 (score_3_x487),
 .score_4 (score_4_x487),
 .score_5 (score_5_x487),
 .score_6 (score_6_x487),
 .score_7 (score_7_x487),
 .score_8 (score_8_x487),
 .score_9 (score_9_x487)
);
 
myram_28X28 #(
.ID(488),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x488),
.W_1(W_1_x488),
.W_2(W_2_x488),
.W_3(W_3_x488),
.W_4(W_4_x488),
.W_5(W_5_x488),
.W_6(W_6_x488),
.W_7(W_7_x488),
.W_8(W_8_x488),
.W_9(W_9_x488)
) u_28X28_x488 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x488),
 .score_0 (score_0_x488),
 .score_1 (score_1_x488),
 .score_2 (score_2_x488),
 .score_3 (score_3_x488),
 .score_4 (score_4_x488),
 .score_5 (score_5_x488),
 .score_6 (score_6_x488),
 .score_7 (score_7_x488),
 .score_8 (score_8_x488),
 .score_9 (score_9_x488)
);
 
myram_28X28 #(
.ID(489),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x489),
.W_1(W_1_x489),
.W_2(W_2_x489),
.W_3(W_3_x489),
.W_4(W_4_x489),
.W_5(W_5_x489),
.W_6(W_6_x489),
.W_7(W_7_x489),
.W_8(W_8_x489),
.W_9(W_9_x489)
) u_28X28_x489 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x489),
 .score_0 (score_0_x489),
 .score_1 (score_1_x489),
 .score_2 (score_2_x489),
 .score_3 (score_3_x489),
 .score_4 (score_4_x489),
 .score_5 (score_5_x489),
 .score_6 (score_6_x489),
 .score_7 (score_7_x489),
 .score_8 (score_8_x489),
 .score_9 (score_9_x489)
);
 
myram_28X28 #(
.ID(490),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x490),
.W_1(W_1_x490),
.W_2(W_2_x490),
.W_3(W_3_x490),
.W_4(W_4_x490),
.W_5(W_5_x490),
.W_6(W_6_x490),
.W_7(W_7_x490),
.W_8(W_8_x490),
.W_9(W_9_x490)
) u_28X28_x490 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x490),
 .score_0 (score_0_x490),
 .score_1 (score_1_x490),
 .score_2 (score_2_x490),
 .score_3 (score_3_x490),
 .score_4 (score_4_x490),
 .score_5 (score_5_x490),
 .score_6 (score_6_x490),
 .score_7 (score_7_x490),
 .score_8 (score_8_x490),
 .score_9 (score_9_x490)
);
 
myram_28X28 #(
.ID(491),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x491),
.W_1(W_1_x491),
.W_2(W_2_x491),
.W_3(W_3_x491),
.W_4(W_4_x491),
.W_5(W_5_x491),
.W_6(W_6_x491),
.W_7(W_7_x491),
.W_8(W_8_x491),
.W_9(W_9_x491)
) u_28X28_x491 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x491),
 .score_0 (score_0_x491),
 .score_1 (score_1_x491),
 .score_2 (score_2_x491),
 .score_3 (score_3_x491),
 .score_4 (score_4_x491),
 .score_5 (score_5_x491),
 .score_6 (score_6_x491),
 .score_7 (score_7_x491),
 .score_8 (score_8_x491),
 .score_9 (score_9_x491)
);
 
myram_28X28 #(
.ID(492),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x492),
.W_1(W_1_x492),
.W_2(W_2_x492),
.W_3(W_3_x492),
.W_4(W_4_x492),
.W_5(W_5_x492),
.W_6(W_6_x492),
.W_7(W_7_x492),
.W_8(W_8_x492),
.W_9(W_9_x492)
) u_28X28_x492 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x492),
 .score_0 (score_0_x492),
 .score_1 (score_1_x492),
 .score_2 (score_2_x492),
 .score_3 (score_3_x492),
 .score_4 (score_4_x492),
 .score_5 (score_5_x492),
 .score_6 (score_6_x492),
 .score_7 (score_7_x492),
 .score_8 (score_8_x492),
 .score_9 (score_9_x492)
);
 
myram_28X28 #(
.ID(493),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x493),
.W_1(W_1_x493),
.W_2(W_2_x493),
.W_3(W_3_x493),
.W_4(W_4_x493),
.W_5(W_5_x493),
.W_6(W_6_x493),
.W_7(W_7_x493),
.W_8(W_8_x493),
.W_9(W_9_x493)
) u_28X28_x493 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x493),
 .score_0 (score_0_x493),
 .score_1 (score_1_x493),
 .score_2 (score_2_x493),
 .score_3 (score_3_x493),
 .score_4 (score_4_x493),
 .score_5 (score_5_x493),
 .score_6 (score_6_x493),
 .score_7 (score_7_x493),
 .score_8 (score_8_x493),
 .score_9 (score_9_x493)
);
 
myram_28X28 #(
.ID(494),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x494),
.W_1(W_1_x494),
.W_2(W_2_x494),
.W_3(W_3_x494),
.W_4(W_4_x494),
.W_5(W_5_x494),
.W_6(W_6_x494),
.W_7(W_7_x494),
.W_8(W_8_x494),
.W_9(W_9_x494)
) u_28X28_x494 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x494),
 .score_0 (score_0_x494),
 .score_1 (score_1_x494),
 .score_2 (score_2_x494),
 .score_3 (score_3_x494),
 .score_4 (score_4_x494),
 .score_5 (score_5_x494),
 .score_6 (score_6_x494),
 .score_7 (score_7_x494),
 .score_8 (score_8_x494),
 .score_9 (score_9_x494)
);
 
myram_28X28 #(
.ID(495),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x495),
.W_1(W_1_x495),
.W_2(W_2_x495),
.W_3(W_3_x495),
.W_4(W_4_x495),
.W_5(W_5_x495),
.W_6(W_6_x495),
.W_7(W_7_x495),
.W_8(W_8_x495),
.W_9(W_9_x495)
) u_28X28_x495 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x495),
 .score_0 (score_0_x495),
 .score_1 (score_1_x495),
 .score_2 (score_2_x495),
 .score_3 (score_3_x495),
 .score_4 (score_4_x495),
 .score_5 (score_5_x495),
 .score_6 (score_6_x495),
 .score_7 (score_7_x495),
 .score_8 (score_8_x495),
 .score_9 (score_9_x495)
);
 
myram_28X28 #(
.ID(496),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x496),
.W_1(W_1_x496),
.W_2(W_2_x496),
.W_3(W_3_x496),
.W_4(W_4_x496),
.W_5(W_5_x496),
.W_6(W_6_x496),
.W_7(W_7_x496),
.W_8(W_8_x496),
.W_9(W_9_x496)
) u_28X28_x496 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x496),
 .score_0 (score_0_x496),
 .score_1 (score_1_x496),
 .score_2 (score_2_x496),
 .score_3 (score_3_x496),
 .score_4 (score_4_x496),
 .score_5 (score_5_x496),
 .score_6 (score_6_x496),
 .score_7 (score_7_x496),
 .score_8 (score_8_x496),
 .score_9 (score_9_x496)
);
 
myram_28X28 #(
.ID(497),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x497),
.W_1(W_1_x497),
.W_2(W_2_x497),
.W_3(W_3_x497),
.W_4(W_4_x497),
.W_5(W_5_x497),
.W_6(W_6_x497),
.W_7(W_7_x497),
.W_8(W_8_x497),
.W_9(W_9_x497)
) u_28X28_x497 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x497),
 .score_0 (score_0_x497),
 .score_1 (score_1_x497),
 .score_2 (score_2_x497),
 .score_3 (score_3_x497),
 .score_4 (score_4_x497),
 .score_5 (score_5_x497),
 .score_6 (score_6_x497),
 .score_7 (score_7_x497),
 .score_8 (score_8_x497),
 .score_9 (score_9_x497)
);
 
myram_28X28 #(
.ID(498),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x498),
.W_1(W_1_x498),
.W_2(W_2_x498),
.W_3(W_3_x498),
.W_4(W_4_x498),
.W_5(W_5_x498),
.W_6(W_6_x498),
.W_7(W_7_x498),
.W_8(W_8_x498),
.W_9(W_9_x498)
) u_28X28_x498 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x498),
 .score_0 (score_0_x498),
 .score_1 (score_1_x498),
 .score_2 (score_2_x498),
 .score_3 (score_3_x498),
 .score_4 (score_4_x498),
 .score_5 (score_5_x498),
 .score_6 (score_6_x498),
 .score_7 (score_7_x498),
 .score_8 (score_8_x498),
 .score_9 (score_9_x498)
);
 
myram_28X28 #(
.ID(499),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x499),
.W_1(W_1_x499),
.W_2(W_2_x499),
.W_3(W_3_x499),
.W_4(W_4_x499),
.W_5(W_5_x499),
.W_6(W_6_x499),
.W_7(W_7_x499),
.W_8(W_8_x499),
.W_9(W_9_x499)
) u_28X28_x499 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x499),
 .score_0 (score_0_x499),
 .score_1 (score_1_x499),
 .score_2 (score_2_x499),
 .score_3 (score_3_x499),
 .score_4 (score_4_x499),
 .score_5 (score_5_x499),
 .score_6 (score_6_x499),
 .score_7 (score_7_x499),
 .score_8 (score_8_x499),
 .score_9 (score_9_x499)
);
 
myram_28X28 #(
.ID(500),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x500),
.W_1(W_1_x500),
.W_2(W_2_x500),
.W_3(W_3_x500),
.W_4(W_4_x500),
.W_5(W_5_x500),
.W_6(W_6_x500),
.W_7(W_7_x500),
.W_8(W_8_x500),
.W_9(W_9_x500)
) u_28X28_x500 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x500),
 .score_0 (score_0_x500),
 .score_1 (score_1_x500),
 .score_2 (score_2_x500),
 .score_3 (score_3_x500),
 .score_4 (score_4_x500),
 .score_5 (score_5_x500),
 .score_6 (score_6_x500),
 .score_7 (score_7_x500),
 .score_8 (score_8_x500),
 .score_9 (score_9_x500)
);
 
myram_28X28 #(
.ID(501),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x501),
.W_1(W_1_x501),
.W_2(W_2_x501),
.W_3(W_3_x501),
.W_4(W_4_x501),
.W_5(W_5_x501),
.W_6(W_6_x501),
.W_7(W_7_x501),
.W_8(W_8_x501),
.W_9(W_9_x501)
) u_28X28_x501 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x501),
 .score_0 (score_0_x501),
 .score_1 (score_1_x501),
 .score_2 (score_2_x501),
 .score_3 (score_3_x501),
 .score_4 (score_4_x501),
 .score_5 (score_5_x501),
 .score_6 (score_6_x501),
 .score_7 (score_7_x501),
 .score_8 (score_8_x501),
 .score_9 (score_9_x501)
);
 
myram_28X28 #(
.ID(502),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x502),
.W_1(W_1_x502),
.W_2(W_2_x502),
.W_3(W_3_x502),
.W_4(W_4_x502),
.W_5(W_5_x502),
.W_6(W_6_x502),
.W_7(W_7_x502),
.W_8(W_8_x502),
.W_9(W_9_x502)
) u_28X28_x502 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x502),
 .score_0 (score_0_x502),
 .score_1 (score_1_x502),
 .score_2 (score_2_x502),
 .score_3 (score_3_x502),
 .score_4 (score_4_x502),
 .score_5 (score_5_x502),
 .score_6 (score_6_x502),
 .score_7 (score_7_x502),
 .score_8 (score_8_x502),
 .score_9 (score_9_x502)
);
 
myram_28X28 #(
.ID(503),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x503),
.W_1(W_1_x503),
.W_2(W_2_x503),
.W_3(W_3_x503),
.W_4(W_4_x503),
.W_5(W_5_x503),
.W_6(W_6_x503),
.W_7(W_7_x503),
.W_8(W_8_x503),
.W_9(W_9_x503)
) u_28X28_x503 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x503),
 .score_0 (score_0_x503),
 .score_1 (score_1_x503),
 .score_2 (score_2_x503),
 .score_3 (score_3_x503),
 .score_4 (score_4_x503),
 .score_5 (score_5_x503),
 .score_6 (score_6_x503),
 .score_7 (score_7_x503),
 .score_8 (score_8_x503),
 .score_9 (score_9_x503)
);
 
myram_28X28 #(
.ID(504),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x504),
.W_1(W_1_x504),
.W_2(W_2_x504),
.W_3(W_3_x504),
.W_4(W_4_x504),
.W_5(W_5_x504),
.W_6(W_6_x504),
.W_7(W_7_x504),
.W_8(W_8_x504),
.W_9(W_9_x504)
) u_28X28_x504 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x504),
 .score_0 (score_0_x504),
 .score_1 (score_1_x504),
 .score_2 (score_2_x504),
 .score_3 (score_3_x504),
 .score_4 (score_4_x504),
 .score_5 (score_5_x504),
 .score_6 (score_6_x504),
 .score_7 (score_7_x504),
 .score_8 (score_8_x504),
 .score_9 (score_9_x504)
);
 
myram_28X28 #(
.ID(505),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x505),
.W_1(W_1_x505),
.W_2(W_2_x505),
.W_3(W_3_x505),
.W_4(W_4_x505),
.W_5(W_5_x505),
.W_6(W_6_x505),
.W_7(W_7_x505),
.W_8(W_8_x505),
.W_9(W_9_x505)
) u_28X28_x505 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x505),
 .score_0 (score_0_x505),
 .score_1 (score_1_x505),
 .score_2 (score_2_x505),
 .score_3 (score_3_x505),
 .score_4 (score_4_x505),
 .score_5 (score_5_x505),
 .score_6 (score_6_x505),
 .score_7 (score_7_x505),
 .score_8 (score_8_x505),
 .score_9 (score_9_x505)
);
 
myram_28X28 #(
.ID(506),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x506),
.W_1(W_1_x506),
.W_2(W_2_x506),
.W_3(W_3_x506),
.W_4(W_4_x506),
.W_5(W_5_x506),
.W_6(W_6_x506),
.W_7(W_7_x506),
.W_8(W_8_x506),
.W_9(W_9_x506)
) u_28X28_x506 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x506),
 .score_0 (score_0_x506),
 .score_1 (score_1_x506),
 .score_2 (score_2_x506),
 .score_3 (score_3_x506),
 .score_4 (score_4_x506),
 .score_5 (score_5_x506),
 .score_6 (score_6_x506),
 .score_7 (score_7_x506),
 .score_8 (score_8_x506),
 .score_9 (score_9_x506)
);
 
myram_28X28 #(
.ID(507),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x507),
.W_1(W_1_x507),
.W_2(W_2_x507),
.W_3(W_3_x507),
.W_4(W_4_x507),
.W_5(W_5_x507),
.W_6(W_6_x507),
.W_7(W_7_x507),
.W_8(W_8_x507),
.W_9(W_9_x507)
) u_28X28_x507 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x507),
 .score_0 (score_0_x507),
 .score_1 (score_1_x507),
 .score_2 (score_2_x507),
 .score_3 (score_3_x507),
 .score_4 (score_4_x507),
 .score_5 (score_5_x507),
 .score_6 (score_6_x507),
 .score_7 (score_7_x507),
 .score_8 (score_8_x507),
 .score_9 (score_9_x507)
);
 
myram_28X28 #(
.ID(508),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x508),
.W_1(W_1_x508),
.W_2(W_2_x508),
.W_3(W_3_x508),
.W_4(W_4_x508),
.W_5(W_5_x508),
.W_6(W_6_x508),
.W_7(W_7_x508),
.W_8(W_8_x508),
.W_9(W_9_x508)
) u_28X28_x508 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x508),
 .score_0 (score_0_x508),
 .score_1 (score_1_x508),
 .score_2 (score_2_x508),
 .score_3 (score_3_x508),
 .score_4 (score_4_x508),
 .score_5 (score_5_x508),
 .score_6 (score_6_x508),
 .score_7 (score_7_x508),
 .score_8 (score_8_x508),
 .score_9 (score_9_x508)
);
 
myram_28X28 #(
.ID(509),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x509),
.W_1(W_1_x509),
.W_2(W_2_x509),
.W_3(W_3_x509),
.W_4(W_4_x509),
.W_5(W_5_x509),
.W_6(W_6_x509),
.W_7(W_7_x509),
.W_8(W_8_x509),
.W_9(W_9_x509)
) u_28X28_x509 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x509),
 .score_0 (score_0_x509),
 .score_1 (score_1_x509),
 .score_2 (score_2_x509),
 .score_3 (score_3_x509),
 .score_4 (score_4_x509),
 .score_5 (score_5_x509),
 .score_6 (score_6_x509),
 .score_7 (score_7_x509),
 .score_8 (score_8_x509),
 .score_9 (score_9_x509)
);
 
myram_28X28 #(
.ID(510),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x510),
.W_1(W_1_x510),
.W_2(W_2_x510),
.W_3(W_3_x510),
.W_4(W_4_x510),
.W_5(W_5_x510),
.W_6(W_6_x510),
.W_7(W_7_x510),
.W_8(W_8_x510),
.W_9(W_9_x510)
) u_28X28_x510 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x510),
 .score_0 (score_0_x510),
 .score_1 (score_1_x510),
 .score_2 (score_2_x510),
 .score_3 (score_3_x510),
 .score_4 (score_4_x510),
 .score_5 (score_5_x510),
 .score_6 (score_6_x510),
 .score_7 (score_7_x510),
 .score_8 (score_8_x510),
 .score_9 (score_9_x510)
);
 
myram_28X28 #(
.ID(511),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x511),
.W_1(W_1_x511),
.W_2(W_2_x511),
.W_3(W_3_x511),
.W_4(W_4_x511),
.W_5(W_5_x511),
.W_6(W_6_x511),
.W_7(W_7_x511),
.W_8(W_8_x511),
.W_9(W_9_x511)
) u_28X28_x511 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x511),
 .score_0 (score_0_x511),
 .score_1 (score_1_x511),
 .score_2 (score_2_x511),
 .score_3 (score_3_x511),
 .score_4 (score_4_x511),
 .score_5 (score_5_x511),
 .score_6 (score_6_x511),
 .score_7 (score_7_x511),
 .score_8 (score_8_x511),
 .score_9 (score_9_x511)
);
 
myram_28X28 #(
.ID(512),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x512),
.W_1(W_1_x512),
.W_2(W_2_x512),
.W_3(W_3_x512),
.W_4(W_4_x512),
.W_5(W_5_x512),
.W_6(W_6_x512),
.W_7(W_7_x512),
.W_8(W_8_x512),
.W_9(W_9_x512)
) u_28X28_x512 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x512),
 .score_0 (score_0_x512),
 .score_1 (score_1_x512),
 .score_2 (score_2_x512),
 .score_3 (score_3_x512),
 .score_4 (score_4_x512),
 .score_5 (score_5_x512),
 .score_6 (score_6_x512),
 .score_7 (score_7_x512),
 .score_8 (score_8_x512),
 .score_9 (score_9_x512)
);
 
myram_28X28 #(
.ID(513),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x513),
.W_1(W_1_x513),
.W_2(W_2_x513),
.W_3(W_3_x513),
.W_4(W_4_x513),
.W_5(W_5_x513),
.W_6(W_6_x513),
.W_7(W_7_x513),
.W_8(W_8_x513),
.W_9(W_9_x513)
) u_28X28_x513 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x513),
 .score_0 (score_0_x513),
 .score_1 (score_1_x513),
 .score_2 (score_2_x513),
 .score_3 (score_3_x513),
 .score_4 (score_4_x513),
 .score_5 (score_5_x513),
 .score_6 (score_6_x513),
 .score_7 (score_7_x513),
 .score_8 (score_8_x513),
 .score_9 (score_9_x513)
);
 
myram_28X28 #(
.ID(514),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x514),
.W_1(W_1_x514),
.W_2(W_2_x514),
.W_3(W_3_x514),
.W_4(W_4_x514),
.W_5(W_5_x514),
.W_6(W_6_x514),
.W_7(W_7_x514),
.W_8(W_8_x514),
.W_9(W_9_x514)
) u_28X28_x514 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x514),
 .score_0 (score_0_x514),
 .score_1 (score_1_x514),
 .score_2 (score_2_x514),
 .score_3 (score_3_x514),
 .score_4 (score_4_x514),
 .score_5 (score_5_x514),
 .score_6 (score_6_x514),
 .score_7 (score_7_x514),
 .score_8 (score_8_x514),
 .score_9 (score_9_x514)
);
 
myram_28X28 #(
.ID(515),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x515),
.W_1(W_1_x515),
.W_2(W_2_x515),
.W_3(W_3_x515),
.W_4(W_4_x515),
.W_5(W_5_x515),
.W_6(W_6_x515),
.W_7(W_7_x515),
.W_8(W_8_x515),
.W_9(W_9_x515)
) u_28X28_x515 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x515),
 .score_0 (score_0_x515),
 .score_1 (score_1_x515),
 .score_2 (score_2_x515),
 .score_3 (score_3_x515),
 .score_4 (score_4_x515),
 .score_5 (score_5_x515),
 .score_6 (score_6_x515),
 .score_7 (score_7_x515),
 .score_8 (score_8_x515),
 .score_9 (score_9_x515)
);
 
myram_28X28 #(
.ID(516),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x516),
.W_1(W_1_x516),
.W_2(W_2_x516),
.W_3(W_3_x516),
.W_4(W_4_x516),
.W_5(W_5_x516),
.W_6(W_6_x516),
.W_7(W_7_x516),
.W_8(W_8_x516),
.W_9(W_9_x516)
) u_28X28_x516 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x516),
 .score_0 (score_0_x516),
 .score_1 (score_1_x516),
 .score_2 (score_2_x516),
 .score_3 (score_3_x516),
 .score_4 (score_4_x516),
 .score_5 (score_5_x516),
 .score_6 (score_6_x516),
 .score_7 (score_7_x516),
 .score_8 (score_8_x516),
 .score_9 (score_9_x516)
);
 
myram_28X28 #(
.ID(517),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x517),
.W_1(W_1_x517),
.W_2(W_2_x517),
.W_3(W_3_x517),
.W_4(W_4_x517),
.W_5(W_5_x517),
.W_6(W_6_x517),
.W_7(W_7_x517),
.W_8(W_8_x517),
.W_9(W_9_x517)
) u_28X28_x517 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x517),
 .score_0 (score_0_x517),
 .score_1 (score_1_x517),
 .score_2 (score_2_x517),
 .score_3 (score_3_x517),
 .score_4 (score_4_x517),
 .score_5 (score_5_x517),
 .score_6 (score_6_x517),
 .score_7 (score_7_x517),
 .score_8 (score_8_x517),
 .score_9 (score_9_x517)
);
 
myram_28X28 #(
.ID(518),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x518),
.W_1(W_1_x518),
.W_2(W_2_x518),
.W_3(W_3_x518),
.W_4(W_4_x518),
.W_5(W_5_x518),
.W_6(W_6_x518),
.W_7(W_7_x518),
.W_8(W_8_x518),
.W_9(W_9_x518)
) u_28X28_x518 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x518),
 .score_0 (score_0_x518),
 .score_1 (score_1_x518),
 .score_2 (score_2_x518),
 .score_3 (score_3_x518),
 .score_4 (score_4_x518),
 .score_5 (score_5_x518),
 .score_6 (score_6_x518),
 .score_7 (score_7_x518),
 .score_8 (score_8_x518),
 .score_9 (score_9_x518)
);
 
myram_28X28 #(
.ID(519),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x519),
.W_1(W_1_x519),
.W_2(W_2_x519),
.W_3(W_3_x519),
.W_4(W_4_x519),
.W_5(W_5_x519),
.W_6(W_6_x519),
.W_7(W_7_x519),
.W_8(W_8_x519),
.W_9(W_9_x519)
) u_28X28_x519 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x519),
 .score_0 (score_0_x519),
 .score_1 (score_1_x519),
 .score_2 (score_2_x519),
 .score_3 (score_3_x519),
 .score_4 (score_4_x519),
 .score_5 (score_5_x519),
 .score_6 (score_6_x519),
 .score_7 (score_7_x519),
 .score_8 (score_8_x519),
 .score_9 (score_9_x519)
);
 
myram_28X28 #(
.ID(520),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x520),
.W_1(W_1_x520),
.W_2(W_2_x520),
.W_3(W_3_x520),
.W_4(W_4_x520),
.W_5(W_5_x520),
.W_6(W_6_x520),
.W_7(W_7_x520),
.W_8(W_8_x520),
.W_9(W_9_x520)
) u_28X28_x520 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x520),
 .score_0 (score_0_x520),
 .score_1 (score_1_x520),
 .score_2 (score_2_x520),
 .score_3 (score_3_x520),
 .score_4 (score_4_x520),
 .score_5 (score_5_x520),
 .score_6 (score_6_x520),
 .score_7 (score_7_x520),
 .score_8 (score_8_x520),
 .score_9 (score_9_x520)
);
 
myram_28X28 #(
.ID(521),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x521),
.W_1(W_1_x521),
.W_2(W_2_x521),
.W_3(W_3_x521),
.W_4(W_4_x521),
.W_5(W_5_x521),
.W_6(W_6_x521),
.W_7(W_7_x521),
.W_8(W_8_x521),
.W_9(W_9_x521)
) u_28X28_x521 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x521),
 .score_0 (score_0_x521),
 .score_1 (score_1_x521),
 .score_2 (score_2_x521),
 .score_3 (score_3_x521),
 .score_4 (score_4_x521),
 .score_5 (score_5_x521),
 .score_6 (score_6_x521),
 .score_7 (score_7_x521),
 .score_8 (score_8_x521),
 .score_9 (score_9_x521)
);
 
myram_28X28 #(
.ID(522),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x522),
.W_1(W_1_x522),
.W_2(W_2_x522),
.W_3(W_3_x522),
.W_4(W_4_x522),
.W_5(W_5_x522),
.W_6(W_6_x522),
.W_7(W_7_x522),
.W_8(W_8_x522),
.W_9(W_9_x522)
) u_28X28_x522 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x522),
 .score_0 (score_0_x522),
 .score_1 (score_1_x522),
 .score_2 (score_2_x522),
 .score_3 (score_3_x522),
 .score_4 (score_4_x522),
 .score_5 (score_5_x522),
 .score_6 (score_6_x522),
 .score_7 (score_7_x522),
 .score_8 (score_8_x522),
 .score_9 (score_9_x522)
);
 
myram_28X28 #(
.ID(523),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x523),
.W_1(W_1_x523),
.W_2(W_2_x523),
.W_3(W_3_x523),
.W_4(W_4_x523),
.W_5(W_5_x523),
.W_6(W_6_x523),
.W_7(W_7_x523),
.W_8(W_8_x523),
.W_9(W_9_x523)
) u_28X28_x523 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x523),
 .score_0 (score_0_x523),
 .score_1 (score_1_x523),
 .score_2 (score_2_x523),
 .score_3 (score_3_x523),
 .score_4 (score_4_x523),
 .score_5 (score_5_x523),
 .score_6 (score_6_x523),
 .score_7 (score_7_x523),
 .score_8 (score_8_x523),
 .score_9 (score_9_x523)
);
 
myram_28X28 #(
.ID(524),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x524),
.W_1(W_1_x524),
.W_2(W_2_x524),
.W_3(W_3_x524),
.W_4(W_4_x524),
.W_5(W_5_x524),
.W_6(W_6_x524),
.W_7(W_7_x524),
.W_8(W_8_x524),
.W_9(W_9_x524)
) u_28X28_x524 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x524),
 .score_0 (score_0_x524),
 .score_1 (score_1_x524),
 .score_2 (score_2_x524),
 .score_3 (score_3_x524),
 .score_4 (score_4_x524),
 .score_5 (score_5_x524),
 .score_6 (score_6_x524),
 .score_7 (score_7_x524),
 .score_8 (score_8_x524),
 .score_9 (score_9_x524)
);
 
myram_28X28 #(
.ID(525),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x525),
.W_1(W_1_x525),
.W_2(W_2_x525),
.W_3(W_3_x525),
.W_4(W_4_x525),
.W_5(W_5_x525),
.W_6(W_6_x525),
.W_7(W_7_x525),
.W_8(W_8_x525),
.W_9(W_9_x525)
) u_28X28_x525 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x525),
 .score_0 (score_0_x525),
 .score_1 (score_1_x525),
 .score_2 (score_2_x525),
 .score_3 (score_3_x525),
 .score_4 (score_4_x525),
 .score_5 (score_5_x525),
 .score_6 (score_6_x525),
 .score_7 (score_7_x525),
 .score_8 (score_8_x525),
 .score_9 (score_9_x525)
);
 
myram_28X28 #(
.ID(526),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x526),
.W_1(W_1_x526),
.W_2(W_2_x526),
.W_3(W_3_x526),
.W_4(W_4_x526),
.W_5(W_5_x526),
.W_6(W_6_x526),
.W_7(W_7_x526),
.W_8(W_8_x526),
.W_9(W_9_x526)
) u_28X28_x526 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x526),
 .score_0 (score_0_x526),
 .score_1 (score_1_x526),
 .score_2 (score_2_x526),
 .score_3 (score_3_x526),
 .score_4 (score_4_x526),
 .score_5 (score_5_x526),
 .score_6 (score_6_x526),
 .score_7 (score_7_x526),
 .score_8 (score_8_x526),
 .score_9 (score_9_x526)
);
 
myram_28X28 #(
.ID(527),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x527),
.W_1(W_1_x527),
.W_2(W_2_x527),
.W_3(W_3_x527),
.W_4(W_4_x527),
.W_5(W_5_x527),
.W_6(W_6_x527),
.W_7(W_7_x527),
.W_8(W_8_x527),
.W_9(W_9_x527)
) u_28X28_x527 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x527),
 .score_0 (score_0_x527),
 .score_1 (score_1_x527),
 .score_2 (score_2_x527),
 .score_3 (score_3_x527),
 .score_4 (score_4_x527),
 .score_5 (score_5_x527),
 .score_6 (score_6_x527),
 .score_7 (score_7_x527),
 .score_8 (score_8_x527),
 .score_9 (score_9_x527)
);
 
myram_28X28 #(
.ID(528),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x528),
.W_1(W_1_x528),
.W_2(W_2_x528),
.W_3(W_3_x528),
.W_4(W_4_x528),
.W_5(W_5_x528),
.W_6(W_6_x528),
.W_7(W_7_x528),
.W_8(W_8_x528),
.W_9(W_9_x528)
) u_28X28_x528 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x528),
 .score_0 (score_0_x528),
 .score_1 (score_1_x528),
 .score_2 (score_2_x528),
 .score_3 (score_3_x528),
 .score_4 (score_4_x528),
 .score_5 (score_5_x528),
 .score_6 (score_6_x528),
 .score_7 (score_7_x528),
 .score_8 (score_8_x528),
 .score_9 (score_9_x528)
);
 
myram_28X28 #(
.ID(529),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x529),
.W_1(W_1_x529),
.W_2(W_2_x529),
.W_3(W_3_x529),
.W_4(W_4_x529),
.W_5(W_5_x529),
.W_6(W_6_x529),
.W_7(W_7_x529),
.W_8(W_8_x529),
.W_9(W_9_x529)
) u_28X28_x529 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x529),
 .score_0 (score_0_x529),
 .score_1 (score_1_x529),
 .score_2 (score_2_x529),
 .score_3 (score_3_x529),
 .score_4 (score_4_x529),
 .score_5 (score_5_x529),
 .score_6 (score_6_x529),
 .score_7 (score_7_x529),
 .score_8 (score_8_x529),
 .score_9 (score_9_x529)
);
 
myram_28X28 #(
.ID(530),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x530),
.W_1(W_1_x530),
.W_2(W_2_x530),
.W_3(W_3_x530),
.W_4(W_4_x530),
.W_5(W_5_x530),
.W_6(W_6_x530),
.W_7(W_7_x530),
.W_8(W_8_x530),
.W_9(W_9_x530)
) u_28X28_x530 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x530),
 .score_0 (score_0_x530),
 .score_1 (score_1_x530),
 .score_2 (score_2_x530),
 .score_3 (score_3_x530),
 .score_4 (score_4_x530),
 .score_5 (score_5_x530),
 .score_6 (score_6_x530),
 .score_7 (score_7_x530),
 .score_8 (score_8_x530),
 .score_9 (score_9_x530)
);
 
myram_28X28 #(
.ID(531),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x531),
.W_1(W_1_x531),
.W_2(W_2_x531),
.W_3(W_3_x531),
.W_4(W_4_x531),
.W_5(W_5_x531),
.W_6(W_6_x531),
.W_7(W_7_x531),
.W_8(W_8_x531),
.W_9(W_9_x531)
) u_28X28_x531 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x531),
 .score_0 (score_0_x531),
 .score_1 (score_1_x531),
 .score_2 (score_2_x531),
 .score_3 (score_3_x531),
 .score_4 (score_4_x531),
 .score_5 (score_5_x531),
 .score_6 (score_6_x531),
 .score_7 (score_7_x531),
 .score_8 (score_8_x531),
 .score_9 (score_9_x531)
);
 
myram_28X28 #(
.ID(532),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x532),
.W_1(W_1_x532),
.W_2(W_2_x532),
.W_3(W_3_x532),
.W_4(W_4_x532),
.W_5(W_5_x532),
.W_6(W_6_x532),
.W_7(W_7_x532),
.W_8(W_8_x532),
.W_9(W_9_x532)
) u_28X28_x532 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x532),
 .score_0 (score_0_x532),
 .score_1 (score_1_x532),
 .score_2 (score_2_x532),
 .score_3 (score_3_x532),
 .score_4 (score_4_x532),
 .score_5 (score_5_x532),
 .score_6 (score_6_x532),
 .score_7 (score_7_x532),
 .score_8 (score_8_x532),
 .score_9 (score_9_x532)
);
 
myram_28X28 #(
.ID(533),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x533),
.W_1(W_1_x533),
.W_2(W_2_x533),
.W_3(W_3_x533),
.W_4(W_4_x533),
.W_5(W_5_x533),
.W_6(W_6_x533),
.W_7(W_7_x533),
.W_8(W_8_x533),
.W_9(W_9_x533)
) u_28X28_x533 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x533),
 .score_0 (score_0_x533),
 .score_1 (score_1_x533),
 .score_2 (score_2_x533),
 .score_3 (score_3_x533),
 .score_4 (score_4_x533),
 .score_5 (score_5_x533),
 .score_6 (score_6_x533),
 .score_7 (score_7_x533),
 .score_8 (score_8_x533),
 .score_9 (score_9_x533)
);
 
myram_28X28 #(
.ID(534),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x534),
.W_1(W_1_x534),
.W_2(W_2_x534),
.W_3(W_3_x534),
.W_4(W_4_x534),
.W_5(W_5_x534),
.W_6(W_6_x534),
.W_7(W_7_x534),
.W_8(W_8_x534),
.W_9(W_9_x534)
) u_28X28_x534 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x534),
 .score_0 (score_0_x534),
 .score_1 (score_1_x534),
 .score_2 (score_2_x534),
 .score_3 (score_3_x534),
 .score_4 (score_4_x534),
 .score_5 (score_5_x534),
 .score_6 (score_6_x534),
 .score_7 (score_7_x534),
 .score_8 (score_8_x534),
 .score_9 (score_9_x534)
);
 
myram_28X28 #(
.ID(535),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x535),
.W_1(W_1_x535),
.W_2(W_2_x535),
.W_3(W_3_x535),
.W_4(W_4_x535),
.W_5(W_5_x535),
.W_6(W_6_x535),
.W_7(W_7_x535),
.W_8(W_8_x535),
.W_9(W_9_x535)
) u_28X28_x535 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x535),
 .score_0 (score_0_x535),
 .score_1 (score_1_x535),
 .score_2 (score_2_x535),
 .score_3 (score_3_x535),
 .score_4 (score_4_x535),
 .score_5 (score_5_x535),
 .score_6 (score_6_x535),
 .score_7 (score_7_x535),
 .score_8 (score_8_x535),
 .score_9 (score_9_x535)
);
 
myram_28X28 #(
.ID(536),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x536),
.W_1(W_1_x536),
.W_2(W_2_x536),
.W_3(W_3_x536),
.W_4(W_4_x536),
.W_5(W_5_x536),
.W_6(W_6_x536),
.W_7(W_7_x536),
.W_8(W_8_x536),
.W_9(W_9_x536)
) u_28X28_x536 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x536),
 .score_0 (score_0_x536),
 .score_1 (score_1_x536),
 .score_2 (score_2_x536),
 .score_3 (score_3_x536),
 .score_4 (score_4_x536),
 .score_5 (score_5_x536),
 .score_6 (score_6_x536),
 .score_7 (score_7_x536),
 .score_8 (score_8_x536),
 .score_9 (score_9_x536)
);
 
myram_28X28 #(
.ID(537),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x537),
.W_1(W_1_x537),
.W_2(W_2_x537),
.W_3(W_3_x537),
.W_4(W_4_x537),
.W_5(W_5_x537),
.W_6(W_6_x537),
.W_7(W_7_x537),
.W_8(W_8_x537),
.W_9(W_9_x537)
) u_28X28_x537 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x537),
 .score_0 (score_0_x537),
 .score_1 (score_1_x537),
 .score_2 (score_2_x537),
 .score_3 (score_3_x537),
 .score_4 (score_4_x537),
 .score_5 (score_5_x537),
 .score_6 (score_6_x537),
 .score_7 (score_7_x537),
 .score_8 (score_8_x537),
 .score_9 (score_9_x537)
);
 
myram_28X28 #(
.ID(538),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x538),
.W_1(W_1_x538),
.W_2(W_2_x538),
.W_3(W_3_x538),
.W_4(W_4_x538),
.W_5(W_5_x538),
.W_6(W_6_x538),
.W_7(W_7_x538),
.W_8(W_8_x538),
.W_9(W_9_x538)
) u_28X28_x538 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x538),
 .score_0 (score_0_x538),
 .score_1 (score_1_x538),
 .score_2 (score_2_x538),
 .score_3 (score_3_x538),
 .score_4 (score_4_x538),
 .score_5 (score_5_x538),
 .score_6 (score_6_x538),
 .score_7 (score_7_x538),
 .score_8 (score_8_x538),
 .score_9 (score_9_x538)
);
 
myram_28X28 #(
.ID(539),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x539),
.W_1(W_1_x539),
.W_2(W_2_x539),
.W_3(W_3_x539),
.W_4(W_4_x539),
.W_5(W_5_x539),
.W_6(W_6_x539),
.W_7(W_7_x539),
.W_8(W_8_x539),
.W_9(W_9_x539)
) u_28X28_x539 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x539),
 .score_0 (score_0_x539),
 .score_1 (score_1_x539),
 .score_2 (score_2_x539),
 .score_3 (score_3_x539),
 .score_4 (score_4_x539),
 .score_5 (score_5_x539),
 .score_6 (score_6_x539),
 .score_7 (score_7_x539),
 .score_8 (score_8_x539),
 .score_9 (score_9_x539)
);
 
myram_28X28 #(
.ID(540),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x540),
.W_1(W_1_x540),
.W_2(W_2_x540),
.W_3(W_3_x540),
.W_4(W_4_x540),
.W_5(W_5_x540),
.W_6(W_6_x540),
.W_7(W_7_x540),
.W_8(W_8_x540),
.W_9(W_9_x540)
) u_28X28_x540 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x540),
 .score_0 (score_0_x540),
 .score_1 (score_1_x540),
 .score_2 (score_2_x540),
 .score_3 (score_3_x540),
 .score_4 (score_4_x540),
 .score_5 (score_5_x540),
 .score_6 (score_6_x540),
 .score_7 (score_7_x540),
 .score_8 (score_8_x540),
 .score_9 (score_9_x540)
);
 
myram_28X28 #(
.ID(541),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x541),
.W_1(W_1_x541),
.W_2(W_2_x541),
.W_3(W_3_x541),
.W_4(W_4_x541),
.W_5(W_5_x541),
.W_6(W_6_x541),
.W_7(W_7_x541),
.W_8(W_8_x541),
.W_9(W_9_x541)
) u_28X28_x541 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x541),
 .score_0 (score_0_x541),
 .score_1 (score_1_x541),
 .score_2 (score_2_x541),
 .score_3 (score_3_x541),
 .score_4 (score_4_x541),
 .score_5 (score_5_x541),
 .score_6 (score_6_x541),
 .score_7 (score_7_x541),
 .score_8 (score_8_x541),
 .score_9 (score_9_x541)
);
 
myram_28X28 #(
.ID(542),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x542),
.W_1(W_1_x542),
.W_2(W_2_x542),
.W_3(W_3_x542),
.W_4(W_4_x542),
.W_5(W_5_x542),
.W_6(W_6_x542),
.W_7(W_7_x542),
.W_8(W_8_x542),
.W_9(W_9_x542)
) u_28X28_x542 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x542),
 .score_0 (score_0_x542),
 .score_1 (score_1_x542),
 .score_2 (score_2_x542),
 .score_3 (score_3_x542),
 .score_4 (score_4_x542),
 .score_5 (score_5_x542),
 .score_6 (score_6_x542),
 .score_7 (score_7_x542),
 .score_8 (score_8_x542),
 .score_9 (score_9_x542)
);
 
myram_28X28 #(
.ID(543),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x543),
.W_1(W_1_x543),
.W_2(W_2_x543),
.W_3(W_3_x543),
.W_4(W_4_x543),
.W_5(W_5_x543),
.W_6(W_6_x543),
.W_7(W_7_x543),
.W_8(W_8_x543),
.W_9(W_9_x543)
) u_28X28_x543 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x543),
 .score_0 (score_0_x543),
 .score_1 (score_1_x543),
 .score_2 (score_2_x543),
 .score_3 (score_3_x543),
 .score_4 (score_4_x543),
 .score_5 (score_5_x543),
 .score_6 (score_6_x543),
 .score_7 (score_7_x543),
 .score_8 (score_8_x543),
 .score_9 (score_9_x543)
);
 
myram_28X28 #(
.ID(544),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x544),
.W_1(W_1_x544),
.W_2(W_2_x544),
.W_3(W_3_x544),
.W_4(W_4_x544),
.W_5(W_5_x544),
.W_6(W_6_x544),
.W_7(W_7_x544),
.W_8(W_8_x544),
.W_9(W_9_x544)
) u_28X28_x544 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x544),
 .score_0 (score_0_x544),
 .score_1 (score_1_x544),
 .score_2 (score_2_x544),
 .score_3 (score_3_x544),
 .score_4 (score_4_x544),
 .score_5 (score_5_x544),
 .score_6 (score_6_x544),
 .score_7 (score_7_x544),
 .score_8 (score_8_x544),
 .score_9 (score_9_x544)
);
 
myram_28X28 #(
.ID(545),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x545),
.W_1(W_1_x545),
.W_2(W_2_x545),
.W_3(W_3_x545),
.W_4(W_4_x545),
.W_5(W_5_x545),
.W_6(W_6_x545),
.W_7(W_7_x545),
.W_8(W_8_x545),
.W_9(W_9_x545)
) u_28X28_x545 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x545),
 .score_0 (score_0_x545),
 .score_1 (score_1_x545),
 .score_2 (score_2_x545),
 .score_3 (score_3_x545),
 .score_4 (score_4_x545),
 .score_5 (score_5_x545),
 .score_6 (score_6_x545),
 .score_7 (score_7_x545),
 .score_8 (score_8_x545),
 .score_9 (score_9_x545)
);
 
myram_28X28 #(
.ID(546),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x546),
.W_1(W_1_x546),
.W_2(W_2_x546),
.W_3(W_3_x546),
.W_4(W_4_x546),
.W_5(W_5_x546),
.W_6(W_6_x546),
.W_7(W_7_x546),
.W_8(W_8_x546),
.W_9(W_9_x546)
) u_28X28_x546 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x546),
 .score_0 (score_0_x546),
 .score_1 (score_1_x546),
 .score_2 (score_2_x546),
 .score_3 (score_3_x546),
 .score_4 (score_4_x546),
 .score_5 (score_5_x546),
 .score_6 (score_6_x546),
 .score_7 (score_7_x546),
 .score_8 (score_8_x546),
 .score_9 (score_9_x546)
);
 
myram_28X28 #(
.ID(547),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x547),
.W_1(W_1_x547),
.W_2(W_2_x547),
.W_3(W_3_x547),
.W_4(W_4_x547),
.W_5(W_5_x547),
.W_6(W_6_x547),
.W_7(W_7_x547),
.W_8(W_8_x547),
.W_9(W_9_x547)
) u_28X28_x547 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x547),
 .score_0 (score_0_x547),
 .score_1 (score_1_x547),
 .score_2 (score_2_x547),
 .score_3 (score_3_x547),
 .score_4 (score_4_x547),
 .score_5 (score_5_x547),
 .score_6 (score_6_x547),
 .score_7 (score_7_x547),
 .score_8 (score_8_x547),
 .score_9 (score_9_x547)
);
 
myram_28X28 #(
.ID(548),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x548),
.W_1(W_1_x548),
.W_2(W_2_x548),
.W_3(W_3_x548),
.W_4(W_4_x548),
.W_5(W_5_x548),
.W_6(W_6_x548),
.W_7(W_7_x548),
.W_8(W_8_x548),
.W_9(W_9_x548)
) u_28X28_x548 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x548),
 .score_0 (score_0_x548),
 .score_1 (score_1_x548),
 .score_2 (score_2_x548),
 .score_3 (score_3_x548),
 .score_4 (score_4_x548),
 .score_5 (score_5_x548),
 .score_6 (score_6_x548),
 .score_7 (score_7_x548),
 .score_8 (score_8_x548),
 .score_9 (score_9_x548)
);
 
myram_28X28 #(
.ID(549),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x549),
.W_1(W_1_x549),
.W_2(W_2_x549),
.W_3(W_3_x549),
.W_4(W_4_x549),
.W_5(W_5_x549),
.W_6(W_6_x549),
.W_7(W_7_x549),
.W_8(W_8_x549),
.W_9(W_9_x549)
) u_28X28_x549 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x549),
 .score_0 (score_0_x549),
 .score_1 (score_1_x549),
 .score_2 (score_2_x549),
 .score_3 (score_3_x549),
 .score_4 (score_4_x549),
 .score_5 (score_5_x549),
 .score_6 (score_6_x549),
 .score_7 (score_7_x549),
 .score_8 (score_8_x549),
 .score_9 (score_9_x549)
);
 
myram_28X28 #(
.ID(550),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x550),
.W_1(W_1_x550),
.W_2(W_2_x550),
.W_3(W_3_x550),
.W_4(W_4_x550),
.W_5(W_5_x550),
.W_6(W_6_x550),
.W_7(W_7_x550),
.W_8(W_8_x550),
.W_9(W_9_x550)
) u_28X28_x550 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x550),
 .score_0 (score_0_x550),
 .score_1 (score_1_x550),
 .score_2 (score_2_x550),
 .score_3 (score_3_x550),
 .score_4 (score_4_x550),
 .score_5 (score_5_x550),
 .score_6 (score_6_x550),
 .score_7 (score_7_x550),
 .score_8 (score_8_x550),
 .score_9 (score_9_x550)
);
 
myram_28X28 #(
.ID(551),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x551),
.W_1(W_1_x551),
.W_2(W_2_x551),
.W_3(W_3_x551),
.W_4(W_4_x551),
.W_5(W_5_x551),
.W_6(W_6_x551),
.W_7(W_7_x551),
.W_8(W_8_x551),
.W_9(W_9_x551)
) u_28X28_x551 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x551),
 .score_0 (score_0_x551),
 .score_1 (score_1_x551),
 .score_2 (score_2_x551),
 .score_3 (score_3_x551),
 .score_4 (score_4_x551),
 .score_5 (score_5_x551),
 .score_6 (score_6_x551),
 .score_7 (score_7_x551),
 .score_8 (score_8_x551),
 .score_9 (score_9_x551)
);
 
myram_28X28 #(
.ID(552),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x552),
.W_1(W_1_x552),
.W_2(W_2_x552),
.W_3(W_3_x552),
.W_4(W_4_x552),
.W_5(W_5_x552),
.W_6(W_6_x552),
.W_7(W_7_x552),
.W_8(W_8_x552),
.W_9(W_9_x552)
) u_28X28_x552 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x552),
 .score_0 (score_0_x552),
 .score_1 (score_1_x552),
 .score_2 (score_2_x552),
 .score_3 (score_3_x552),
 .score_4 (score_4_x552),
 .score_5 (score_5_x552),
 .score_6 (score_6_x552),
 .score_7 (score_7_x552),
 .score_8 (score_8_x552),
 .score_9 (score_9_x552)
);
 
myram_28X28 #(
.ID(553),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x553),
.W_1(W_1_x553),
.W_2(W_2_x553),
.W_3(W_3_x553),
.W_4(W_4_x553),
.W_5(W_5_x553),
.W_6(W_6_x553),
.W_7(W_7_x553),
.W_8(W_8_x553),
.W_9(W_9_x553)
) u_28X28_x553 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x553),
 .score_0 (score_0_x553),
 .score_1 (score_1_x553),
 .score_2 (score_2_x553),
 .score_3 (score_3_x553),
 .score_4 (score_4_x553),
 .score_5 (score_5_x553),
 .score_6 (score_6_x553),
 .score_7 (score_7_x553),
 .score_8 (score_8_x553),
 .score_9 (score_9_x553)
);
 
myram_28X28 #(
.ID(554),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x554),
.W_1(W_1_x554),
.W_2(W_2_x554),
.W_3(W_3_x554),
.W_4(W_4_x554),
.W_5(W_5_x554),
.W_6(W_6_x554),
.W_7(W_7_x554),
.W_8(W_8_x554),
.W_9(W_9_x554)
) u_28X28_x554 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x554),
 .score_0 (score_0_x554),
 .score_1 (score_1_x554),
 .score_2 (score_2_x554),
 .score_3 (score_3_x554),
 .score_4 (score_4_x554),
 .score_5 (score_5_x554),
 .score_6 (score_6_x554),
 .score_7 (score_7_x554),
 .score_8 (score_8_x554),
 .score_9 (score_9_x554)
);
 
myram_28X28 #(
.ID(555),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x555),
.W_1(W_1_x555),
.W_2(W_2_x555),
.W_3(W_3_x555),
.W_4(W_4_x555),
.W_5(W_5_x555),
.W_6(W_6_x555),
.W_7(W_7_x555),
.W_8(W_8_x555),
.W_9(W_9_x555)
) u_28X28_x555 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x555),
 .score_0 (score_0_x555),
 .score_1 (score_1_x555),
 .score_2 (score_2_x555),
 .score_3 (score_3_x555),
 .score_4 (score_4_x555),
 .score_5 (score_5_x555),
 .score_6 (score_6_x555),
 .score_7 (score_7_x555),
 .score_8 (score_8_x555),
 .score_9 (score_9_x555)
);
 
myram_28X28 #(
.ID(556),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x556),
.W_1(W_1_x556),
.W_2(W_2_x556),
.W_3(W_3_x556),
.W_4(W_4_x556),
.W_5(W_5_x556),
.W_6(W_6_x556),
.W_7(W_7_x556),
.W_8(W_8_x556),
.W_9(W_9_x556)
) u_28X28_x556 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x556),
 .score_0 (score_0_x556),
 .score_1 (score_1_x556),
 .score_2 (score_2_x556),
 .score_3 (score_3_x556),
 .score_4 (score_4_x556),
 .score_5 (score_5_x556),
 .score_6 (score_6_x556),
 .score_7 (score_7_x556),
 .score_8 (score_8_x556),
 .score_9 (score_9_x556)
);
 
myram_28X28 #(
.ID(557),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x557),
.W_1(W_1_x557),
.W_2(W_2_x557),
.W_3(W_3_x557),
.W_4(W_4_x557),
.W_5(W_5_x557),
.W_6(W_6_x557),
.W_7(W_7_x557),
.W_8(W_8_x557),
.W_9(W_9_x557)
) u_28X28_x557 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x557),
 .score_0 (score_0_x557),
 .score_1 (score_1_x557),
 .score_2 (score_2_x557),
 .score_3 (score_3_x557),
 .score_4 (score_4_x557),
 .score_5 (score_5_x557),
 .score_6 (score_6_x557),
 .score_7 (score_7_x557),
 .score_8 (score_8_x557),
 .score_9 (score_9_x557)
);
 
myram_28X28 #(
.ID(558),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x558),
.W_1(W_1_x558),
.W_2(W_2_x558),
.W_3(W_3_x558),
.W_4(W_4_x558),
.W_5(W_5_x558),
.W_6(W_6_x558),
.W_7(W_7_x558),
.W_8(W_8_x558),
.W_9(W_9_x558)
) u_28X28_x558 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x558),
 .score_0 (score_0_x558),
 .score_1 (score_1_x558),
 .score_2 (score_2_x558),
 .score_3 (score_3_x558),
 .score_4 (score_4_x558),
 .score_5 (score_5_x558),
 .score_6 (score_6_x558),
 .score_7 (score_7_x558),
 .score_8 (score_8_x558),
 .score_9 (score_9_x558)
);
 
myram_28X28 #(
.ID(559),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x559),
.W_1(W_1_x559),
.W_2(W_2_x559),
.W_3(W_3_x559),
.W_4(W_4_x559),
.W_5(W_5_x559),
.W_6(W_6_x559),
.W_7(W_7_x559),
.W_8(W_8_x559),
.W_9(W_9_x559)
) u_28X28_x559 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x559),
 .score_0 (score_0_x559),
 .score_1 (score_1_x559),
 .score_2 (score_2_x559),
 .score_3 (score_3_x559),
 .score_4 (score_4_x559),
 .score_5 (score_5_x559),
 .score_6 (score_6_x559),
 .score_7 (score_7_x559),
 .score_8 (score_8_x559),
 .score_9 (score_9_x559)
);
 
myram_28X28 #(
.ID(560),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x560),
.W_1(W_1_x560),
.W_2(W_2_x560),
.W_3(W_3_x560),
.W_4(W_4_x560),
.W_5(W_5_x560),
.W_6(W_6_x560),
.W_7(W_7_x560),
.W_8(W_8_x560),
.W_9(W_9_x560)
) u_28X28_x560 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x560),
 .score_0 (score_0_x560),
 .score_1 (score_1_x560),
 .score_2 (score_2_x560),
 .score_3 (score_3_x560),
 .score_4 (score_4_x560),
 .score_5 (score_5_x560),
 .score_6 (score_6_x560),
 .score_7 (score_7_x560),
 .score_8 (score_8_x560),
 .score_9 (score_9_x560)
);
 
myram_28X28 #(
.ID(561),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x561),
.W_1(W_1_x561),
.W_2(W_2_x561),
.W_3(W_3_x561),
.W_4(W_4_x561),
.W_5(W_5_x561),
.W_6(W_6_x561),
.W_7(W_7_x561),
.W_8(W_8_x561),
.W_9(W_9_x561)
) u_28X28_x561 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x561),
 .score_0 (score_0_x561),
 .score_1 (score_1_x561),
 .score_2 (score_2_x561),
 .score_3 (score_3_x561),
 .score_4 (score_4_x561),
 .score_5 (score_5_x561),
 .score_6 (score_6_x561),
 .score_7 (score_7_x561),
 .score_8 (score_8_x561),
 .score_9 (score_9_x561)
);
 
myram_28X28 #(
.ID(562),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x562),
.W_1(W_1_x562),
.W_2(W_2_x562),
.W_3(W_3_x562),
.W_4(W_4_x562),
.W_5(W_5_x562),
.W_6(W_6_x562),
.W_7(W_7_x562),
.W_8(W_8_x562),
.W_9(W_9_x562)
) u_28X28_x562 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x562),
 .score_0 (score_0_x562),
 .score_1 (score_1_x562),
 .score_2 (score_2_x562),
 .score_3 (score_3_x562),
 .score_4 (score_4_x562),
 .score_5 (score_5_x562),
 .score_6 (score_6_x562),
 .score_7 (score_7_x562),
 .score_8 (score_8_x562),
 .score_9 (score_9_x562)
);
 
myram_28X28 #(
.ID(563),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x563),
.W_1(W_1_x563),
.W_2(W_2_x563),
.W_3(W_3_x563),
.W_4(W_4_x563),
.W_5(W_5_x563),
.W_6(W_6_x563),
.W_7(W_7_x563),
.W_8(W_8_x563),
.W_9(W_9_x563)
) u_28X28_x563 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x563),
 .score_0 (score_0_x563),
 .score_1 (score_1_x563),
 .score_2 (score_2_x563),
 .score_3 (score_3_x563),
 .score_4 (score_4_x563),
 .score_5 (score_5_x563),
 .score_6 (score_6_x563),
 .score_7 (score_7_x563),
 .score_8 (score_8_x563),
 .score_9 (score_9_x563)
);
 
myram_28X28 #(
.ID(564),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x564),
.W_1(W_1_x564),
.W_2(W_2_x564),
.W_3(W_3_x564),
.W_4(W_4_x564),
.W_5(W_5_x564),
.W_6(W_6_x564),
.W_7(W_7_x564),
.W_8(W_8_x564),
.W_9(W_9_x564)
) u_28X28_x564 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x564),
 .score_0 (score_0_x564),
 .score_1 (score_1_x564),
 .score_2 (score_2_x564),
 .score_3 (score_3_x564),
 .score_4 (score_4_x564),
 .score_5 (score_5_x564),
 .score_6 (score_6_x564),
 .score_7 (score_7_x564),
 .score_8 (score_8_x564),
 .score_9 (score_9_x564)
);
 
myram_28X28 #(
.ID(565),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x565),
.W_1(W_1_x565),
.W_2(W_2_x565),
.W_3(W_3_x565),
.W_4(W_4_x565),
.W_5(W_5_x565),
.W_6(W_6_x565),
.W_7(W_7_x565),
.W_8(W_8_x565),
.W_9(W_9_x565)
) u_28X28_x565 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x565),
 .score_0 (score_0_x565),
 .score_1 (score_1_x565),
 .score_2 (score_2_x565),
 .score_3 (score_3_x565),
 .score_4 (score_4_x565),
 .score_5 (score_5_x565),
 .score_6 (score_6_x565),
 .score_7 (score_7_x565),
 .score_8 (score_8_x565),
 .score_9 (score_9_x565)
);
 
myram_28X28 #(
.ID(566),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x566),
.W_1(W_1_x566),
.W_2(W_2_x566),
.W_3(W_3_x566),
.W_4(W_4_x566),
.W_5(W_5_x566),
.W_6(W_6_x566),
.W_7(W_7_x566),
.W_8(W_8_x566),
.W_9(W_9_x566)
) u_28X28_x566 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x566),
 .score_0 (score_0_x566),
 .score_1 (score_1_x566),
 .score_2 (score_2_x566),
 .score_3 (score_3_x566),
 .score_4 (score_4_x566),
 .score_5 (score_5_x566),
 .score_6 (score_6_x566),
 .score_7 (score_7_x566),
 .score_8 (score_8_x566),
 .score_9 (score_9_x566)
);
 
myram_28X28 #(
.ID(567),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x567),
.W_1(W_1_x567),
.W_2(W_2_x567),
.W_3(W_3_x567),
.W_4(W_4_x567),
.W_5(W_5_x567),
.W_6(W_6_x567),
.W_7(W_7_x567),
.W_8(W_8_x567),
.W_9(W_9_x567)
) u_28X28_x567 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x567),
 .score_0 (score_0_x567),
 .score_1 (score_1_x567),
 .score_2 (score_2_x567),
 .score_3 (score_3_x567),
 .score_4 (score_4_x567),
 .score_5 (score_5_x567),
 .score_6 (score_6_x567),
 .score_7 (score_7_x567),
 .score_8 (score_8_x567),
 .score_9 (score_9_x567)
);
 
myram_28X28 #(
.ID(568),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x568),
.W_1(W_1_x568),
.W_2(W_2_x568),
.W_3(W_3_x568),
.W_4(W_4_x568),
.W_5(W_5_x568),
.W_6(W_6_x568),
.W_7(W_7_x568),
.W_8(W_8_x568),
.W_9(W_9_x568)
) u_28X28_x568 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x568),
 .score_0 (score_0_x568),
 .score_1 (score_1_x568),
 .score_2 (score_2_x568),
 .score_3 (score_3_x568),
 .score_4 (score_4_x568),
 .score_5 (score_5_x568),
 .score_6 (score_6_x568),
 .score_7 (score_7_x568),
 .score_8 (score_8_x568),
 .score_9 (score_9_x568)
);
 
myram_28X28 #(
.ID(569),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x569),
.W_1(W_1_x569),
.W_2(W_2_x569),
.W_3(W_3_x569),
.W_4(W_4_x569),
.W_5(W_5_x569),
.W_6(W_6_x569),
.W_7(W_7_x569),
.W_8(W_8_x569),
.W_9(W_9_x569)
) u_28X28_x569 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x569),
 .score_0 (score_0_x569),
 .score_1 (score_1_x569),
 .score_2 (score_2_x569),
 .score_3 (score_3_x569),
 .score_4 (score_4_x569),
 .score_5 (score_5_x569),
 .score_6 (score_6_x569),
 .score_7 (score_7_x569),
 .score_8 (score_8_x569),
 .score_9 (score_9_x569)
);
 
myram_28X28 #(
.ID(570),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x570),
.W_1(W_1_x570),
.W_2(W_2_x570),
.W_3(W_3_x570),
.W_4(W_4_x570),
.W_5(W_5_x570),
.W_6(W_6_x570),
.W_7(W_7_x570),
.W_8(W_8_x570),
.W_9(W_9_x570)
) u_28X28_x570 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x570),
 .score_0 (score_0_x570),
 .score_1 (score_1_x570),
 .score_2 (score_2_x570),
 .score_3 (score_3_x570),
 .score_4 (score_4_x570),
 .score_5 (score_5_x570),
 .score_6 (score_6_x570),
 .score_7 (score_7_x570),
 .score_8 (score_8_x570),
 .score_9 (score_9_x570)
);
 
myram_28X28 #(
.ID(571),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x571),
.W_1(W_1_x571),
.W_2(W_2_x571),
.W_3(W_3_x571),
.W_4(W_4_x571),
.W_5(W_5_x571),
.W_6(W_6_x571),
.W_7(W_7_x571),
.W_8(W_8_x571),
.W_9(W_9_x571)
) u_28X28_x571 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x571),
 .score_0 (score_0_x571),
 .score_1 (score_1_x571),
 .score_2 (score_2_x571),
 .score_3 (score_3_x571),
 .score_4 (score_4_x571),
 .score_5 (score_5_x571),
 .score_6 (score_6_x571),
 .score_7 (score_7_x571),
 .score_8 (score_8_x571),
 .score_9 (score_9_x571)
);
 
myram_28X28 #(
.ID(572),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x572),
.W_1(W_1_x572),
.W_2(W_2_x572),
.W_3(W_3_x572),
.W_4(W_4_x572),
.W_5(W_5_x572),
.W_6(W_6_x572),
.W_7(W_7_x572),
.W_8(W_8_x572),
.W_9(W_9_x572)
) u_28X28_x572 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x572),
 .score_0 (score_0_x572),
 .score_1 (score_1_x572),
 .score_2 (score_2_x572),
 .score_3 (score_3_x572),
 .score_4 (score_4_x572),
 .score_5 (score_5_x572),
 .score_6 (score_6_x572),
 .score_7 (score_7_x572),
 .score_8 (score_8_x572),
 .score_9 (score_9_x572)
);
 
myram_28X28 #(
.ID(573),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x573),
.W_1(W_1_x573),
.W_2(W_2_x573),
.W_3(W_3_x573),
.W_4(W_4_x573),
.W_5(W_5_x573),
.W_6(W_6_x573),
.W_7(W_7_x573),
.W_8(W_8_x573),
.W_9(W_9_x573)
) u_28X28_x573 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x573),
 .score_0 (score_0_x573),
 .score_1 (score_1_x573),
 .score_2 (score_2_x573),
 .score_3 (score_3_x573),
 .score_4 (score_4_x573),
 .score_5 (score_5_x573),
 .score_6 (score_6_x573),
 .score_7 (score_7_x573),
 .score_8 (score_8_x573),
 .score_9 (score_9_x573)
);
 
myram_28X28 #(
.ID(574),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x574),
.W_1(W_1_x574),
.W_2(W_2_x574),
.W_3(W_3_x574),
.W_4(W_4_x574),
.W_5(W_5_x574),
.W_6(W_6_x574),
.W_7(W_7_x574),
.W_8(W_8_x574),
.W_9(W_9_x574)
) u_28X28_x574 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x574),
 .score_0 (score_0_x574),
 .score_1 (score_1_x574),
 .score_2 (score_2_x574),
 .score_3 (score_3_x574),
 .score_4 (score_4_x574),
 .score_5 (score_5_x574),
 .score_6 (score_6_x574),
 .score_7 (score_7_x574),
 .score_8 (score_8_x574),
 .score_9 (score_9_x574)
);
 
myram_28X28 #(
.ID(575),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x575),
.W_1(W_1_x575),
.W_2(W_2_x575),
.W_3(W_3_x575),
.W_4(W_4_x575),
.W_5(W_5_x575),
.W_6(W_6_x575),
.W_7(W_7_x575),
.W_8(W_8_x575),
.W_9(W_9_x575)
) u_28X28_x575 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x575),
 .score_0 (score_0_x575),
 .score_1 (score_1_x575),
 .score_2 (score_2_x575),
 .score_3 (score_3_x575),
 .score_4 (score_4_x575),
 .score_5 (score_5_x575),
 .score_6 (score_6_x575),
 .score_7 (score_7_x575),
 .score_8 (score_8_x575),
 .score_9 (score_9_x575)
);
 
myram_28X28 #(
.ID(576),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x576),
.W_1(W_1_x576),
.W_2(W_2_x576),
.W_3(W_3_x576),
.W_4(W_4_x576),
.W_5(W_5_x576),
.W_6(W_6_x576),
.W_7(W_7_x576),
.W_8(W_8_x576),
.W_9(W_9_x576)
) u_28X28_x576 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x576),
 .score_0 (score_0_x576),
 .score_1 (score_1_x576),
 .score_2 (score_2_x576),
 .score_3 (score_3_x576),
 .score_4 (score_4_x576),
 .score_5 (score_5_x576),
 .score_6 (score_6_x576),
 .score_7 (score_7_x576),
 .score_8 (score_8_x576),
 .score_9 (score_9_x576)
);
 
myram_28X28 #(
.ID(577),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x577),
.W_1(W_1_x577),
.W_2(W_2_x577),
.W_3(W_3_x577),
.W_4(W_4_x577),
.W_5(W_5_x577),
.W_6(W_6_x577),
.W_7(W_7_x577),
.W_8(W_8_x577),
.W_9(W_9_x577)
) u_28X28_x577 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x577),
 .score_0 (score_0_x577),
 .score_1 (score_1_x577),
 .score_2 (score_2_x577),
 .score_3 (score_3_x577),
 .score_4 (score_4_x577),
 .score_5 (score_5_x577),
 .score_6 (score_6_x577),
 .score_7 (score_7_x577),
 .score_8 (score_8_x577),
 .score_9 (score_9_x577)
);
 
myram_28X28 #(
.ID(578),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x578),
.W_1(W_1_x578),
.W_2(W_2_x578),
.W_3(W_3_x578),
.W_4(W_4_x578),
.W_5(W_5_x578),
.W_6(W_6_x578),
.W_7(W_7_x578),
.W_8(W_8_x578),
.W_9(W_9_x578)
) u_28X28_x578 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x578),
 .score_0 (score_0_x578),
 .score_1 (score_1_x578),
 .score_2 (score_2_x578),
 .score_3 (score_3_x578),
 .score_4 (score_4_x578),
 .score_5 (score_5_x578),
 .score_6 (score_6_x578),
 .score_7 (score_7_x578),
 .score_8 (score_8_x578),
 .score_9 (score_9_x578)
);
 
myram_28X28 #(
.ID(579),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x579),
.W_1(W_1_x579),
.W_2(W_2_x579),
.W_3(W_3_x579),
.W_4(W_4_x579),
.W_5(W_5_x579),
.W_6(W_6_x579),
.W_7(W_7_x579),
.W_8(W_8_x579),
.W_9(W_9_x579)
) u_28X28_x579 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x579),
 .score_0 (score_0_x579),
 .score_1 (score_1_x579),
 .score_2 (score_2_x579),
 .score_3 (score_3_x579),
 .score_4 (score_4_x579),
 .score_5 (score_5_x579),
 .score_6 (score_6_x579),
 .score_7 (score_7_x579),
 .score_8 (score_8_x579),
 .score_9 (score_9_x579)
);
 
myram_28X28 #(
.ID(580),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x580),
.W_1(W_1_x580),
.W_2(W_2_x580),
.W_3(W_3_x580),
.W_4(W_4_x580),
.W_5(W_5_x580),
.W_6(W_6_x580),
.W_7(W_7_x580),
.W_8(W_8_x580),
.W_9(W_9_x580)
) u_28X28_x580 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x580),
 .score_0 (score_0_x580),
 .score_1 (score_1_x580),
 .score_2 (score_2_x580),
 .score_3 (score_3_x580),
 .score_4 (score_4_x580),
 .score_5 (score_5_x580),
 .score_6 (score_6_x580),
 .score_7 (score_7_x580),
 .score_8 (score_8_x580),
 .score_9 (score_9_x580)
);
 
myram_28X28 #(
.ID(581),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x581),
.W_1(W_1_x581),
.W_2(W_2_x581),
.W_3(W_3_x581),
.W_4(W_4_x581),
.W_5(W_5_x581),
.W_6(W_6_x581),
.W_7(W_7_x581),
.W_8(W_8_x581),
.W_9(W_9_x581)
) u_28X28_x581 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x581),
 .score_0 (score_0_x581),
 .score_1 (score_1_x581),
 .score_2 (score_2_x581),
 .score_3 (score_3_x581),
 .score_4 (score_4_x581),
 .score_5 (score_5_x581),
 .score_6 (score_6_x581),
 .score_7 (score_7_x581),
 .score_8 (score_8_x581),
 .score_9 (score_9_x581)
);
 
myram_28X28 #(
.ID(582),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x582),
.W_1(W_1_x582),
.W_2(W_2_x582),
.W_3(W_3_x582),
.W_4(W_4_x582),
.W_5(W_5_x582),
.W_6(W_6_x582),
.W_7(W_7_x582),
.W_8(W_8_x582),
.W_9(W_9_x582)
) u_28X28_x582 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x582),
 .score_0 (score_0_x582),
 .score_1 (score_1_x582),
 .score_2 (score_2_x582),
 .score_3 (score_3_x582),
 .score_4 (score_4_x582),
 .score_5 (score_5_x582),
 .score_6 (score_6_x582),
 .score_7 (score_7_x582),
 .score_8 (score_8_x582),
 .score_9 (score_9_x582)
);
 
myram_28X28 #(
.ID(583),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x583),
.W_1(W_1_x583),
.W_2(W_2_x583),
.W_3(W_3_x583),
.W_4(W_4_x583),
.W_5(W_5_x583),
.W_6(W_6_x583),
.W_7(W_7_x583),
.W_8(W_8_x583),
.W_9(W_9_x583)
) u_28X28_x583 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x583),
 .score_0 (score_0_x583),
 .score_1 (score_1_x583),
 .score_2 (score_2_x583),
 .score_3 (score_3_x583),
 .score_4 (score_4_x583),
 .score_5 (score_5_x583),
 .score_6 (score_6_x583),
 .score_7 (score_7_x583),
 .score_8 (score_8_x583),
 .score_9 (score_9_x583)
);
 
myram_28X28 #(
.ID(584),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x584),
.W_1(W_1_x584),
.W_2(W_2_x584),
.W_3(W_3_x584),
.W_4(W_4_x584),
.W_5(W_5_x584),
.W_6(W_6_x584),
.W_7(W_7_x584),
.W_8(W_8_x584),
.W_9(W_9_x584)
) u_28X28_x584 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x584),
 .score_0 (score_0_x584),
 .score_1 (score_1_x584),
 .score_2 (score_2_x584),
 .score_3 (score_3_x584),
 .score_4 (score_4_x584),
 .score_5 (score_5_x584),
 .score_6 (score_6_x584),
 .score_7 (score_7_x584),
 .score_8 (score_8_x584),
 .score_9 (score_9_x584)
);
 
myram_28X28 #(
.ID(585),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x585),
.W_1(W_1_x585),
.W_2(W_2_x585),
.W_3(W_3_x585),
.W_4(W_4_x585),
.W_5(W_5_x585),
.W_6(W_6_x585),
.W_7(W_7_x585),
.W_8(W_8_x585),
.W_9(W_9_x585)
) u_28X28_x585 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x585),
 .score_0 (score_0_x585),
 .score_1 (score_1_x585),
 .score_2 (score_2_x585),
 .score_3 (score_3_x585),
 .score_4 (score_4_x585),
 .score_5 (score_5_x585),
 .score_6 (score_6_x585),
 .score_7 (score_7_x585),
 .score_8 (score_8_x585),
 .score_9 (score_9_x585)
);
 
myram_28X28 #(
.ID(586),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x586),
.W_1(W_1_x586),
.W_2(W_2_x586),
.W_3(W_3_x586),
.W_4(W_4_x586),
.W_5(W_5_x586),
.W_6(W_6_x586),
.W_7(W_7_x586),
.W_8(W_8_x586),
.W_9(W_9_x586)
) u_28X28_x586 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x586),
 .score_0 (score_0_x586),
 .score_1 (score_1_x586),
 .score_2 (score_2_x586),
 .score_3 (score_3_x586),
 .score_4 (score_4_x586),
 .score_5 (score_5_x586),
 .score_6 (score_6_x586),
 .score_7 (score_7_x586),
 .score_8 (score_8_x586),
 .score_9 (score_9_x586)
);
 
myram_28X28 #(
.ID(587),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x587),
.W_1(W_1_x587),
.W_2(W_2_x587),
.W_3(W_3_x587),
.W_4(W_4_x587),
.W_5(W_5_x587),
.W_6(W_6_x587),
.W_7(W_7_x587),
.W_8(W_8_x587),
.W_9(W_9_x587)
) u_28X28_x587 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x587),
 .score_0 (score_0_x587),
 .score_1 (score_1_x587),
 .score_2 (score_2_x587),
 .score_3 (score_3_x587),
 .score_4 (score_4_x587),
 .score_5 (score_5_x587),
 .score_6 (score_6_x587),
 .score_7 (score_7_x587),
 .score_8 (score_8_x587),
 .score_9 (score_9_x587)
);
 
myram_28X28 #(
.ID(588),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x588),
.W_1(W_1_x588),
.W_2(W_2_x588),
.W_3(W_3_x588),
.W_4(W_4_x588),
.W_5(W_5_x588),
.W_6(W_6_x588),
.W_7(W_7_x588),
.W_8(W_8_x588),
.W_9(W_9_x588)
) u_28X28_x588 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x588),
 .score_0 (score_0_x588),
 .score_1 (score_1_x588),
 .score_2 (score_2_x588),
 .score_3 (score_3_x588),
 .score_4 (score_4_x588),
 .score_5 (score_5_x588),
 .score_6 (score_6_x588),
 .score_7 (score_7_x588),
 .score_8 (score_8_x588),
 .score_9 (score_9_x588)
);
 
myram_28X28 #(
.ID(589),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x589),
.W_1(W_1_x589),
.W_2(W_2_x589),
.W_3(W_3_x589),
.W_4(W_4_x589),
.W_5(W_5_x589),
.W_6(W_6_x589),
.W_7(W_7_x589),
.W_8(W_8_x589),
.W_9(W_9_x589)
) u_28X28_x589 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x589),
 .score_0 (score_0_x589),
 .score_1 (score_1_x589),
 .score_2 (score_2_x589),
 .score_3 (score_3_x589),
 .score_4 (score_4_x589),
 .score_5 (score_5_x589),
 .score_6 (score_6_x589),
 .score_7 (score_7_x589),
 .score_8 (score_8_x589),
 .score_9 (score_9_x589)
);
 
myram_28X28 #(
.ID(590),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x590),
.W_1(W_1_x590),
.W_2(W_2_x590),
.W_3(W_3_x590),
.W_4(W_4_x590),
.W_5(W_5_x590),
.W_6(W_6_x590),
.W_7(W_7_x590),
.W_8(W_8_x590),
.W_9(W_9_x590)
) u_28X28_x590 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x590),
 .score_0 (score_0_x590),
 .score_1 (score_1_x590),
 .score_2 (score_2_x590),
 .score_3 (score_3_x590),
 .score_4 (score_4_x590),
 .score_5 (score_5_x590),
 .score_6 (score_6_x590),
 .score_7 (score_7_x590),
 .score_8 (score_8_x590),
 .score_9 (score_9_x590)
);
 
myram_28X28 #(
.ID(591),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x591),
.W_1(W_1_x591),
.W_2(W_2_x591),
.W_3(W_3_x591),
.W_4(W_4_x591),
.W_5(W_5_x591),
.W_6(W_6_x591),
.W_7(W_7_x591),
.W_8(W_8_x591),
.W_9(W_9_x591)
) u_28X28_x591 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x591),
 .score_0 (score_0_x591),
 .score_1 (score_1_x591),
 .score_2 (score_2_x591),
 .score_3 (score_3_x591),
 .score_4 (score_4_x591),
 .score_5 (score_5_x591),
 .score_6 (score_6_x591),
 .score_7 (score_7_x591),
 .score_8 (score_8_x591),
 .score_9 (score_9_x591)
);
 
myram_28X28 #(
.ID(592),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x592),
.W_1(W_1_x592),
.W_2(W_2_x592),
.W_3(W_3_x592),
.W_4(W_4_x592),
.W_5(W_5_x592),
.W_6(W_6_x592),
.W_7(W_7_x592),
.W_8(W_8_x592),
.W_9(W_9_x592)
) u_28X28_x592 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x592),
 .score_0 (score_0_x592),
 .score_1 (score_1_x592),
 .score_2 (score_2_x592),
 .score_3 (score_3_x592),
 .score_4 (score_4_x592),
 .score_5 (score_5_x592),
 .score_6 (score_6_x592),
 .score_7 (score_7_x592),
 .score_8 (score_8_x592),
 .score_9 (score_9_x592)
);
 
myram_28X28 #(
.ID(593),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x593),
.W_1(W_1_x593),
.W_2(W_2_x593),
.W_3(W_3_x593),
.W_4(W_4_x593),
.W_5(W_5_x593),
.W_6(W_6_x593),
.W_7(W_7_x593),
.W_8(W_8_x593),
.W_9(W_9_x593)
) u_28X28_x593 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x593),
 .score_0 (score_0_x593),
 .score_1 (score_1_x593),
 .score_2 (score_2_x593),
 .score_3 (score_3_x593),
 .score_4 (score_4_x593),
 .score_5 (score_5_x593),
 .score_6 (score_6_x593),
 .score_7 (score_7_x593),
 .score_8 (score_8_x593),
 .score_9 (score_9_x593)
);
 
myram_28X28 #(
.ID(594),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x594),
.W_1(W_1_x594),
.W_2(W_2_x594),
.W_3(W_3_x594),
.W_4(W_4_x594),
.W_5(W_5_x594),
.W_6(W_6_x594),
.W_7(W_7_x594),
.W_8(W_8_x594),
.W_9(W_9_x594)
) u_28X28_x594 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x594),
 .score_0 (score_0_x594),
 .score_1 (score_1_x594),
 .score_2 (score_2_x594),
 .score_3 (score_3_x594),
 .score_4 (score_4_x594),
 .score_5 (score_5_x594),
 .score_6 (score_6_x594),
 .score_7 (score_7_x594),
 .score_8 (score_8_x594),
 .score_9 (score_9_x594)
);
 
myram_28X28 #(
.ID(595),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x595),
.W_1(W_1_x595),
.W_2(W_2_x595),
.W_3(W_3_x595),
.W_4(W_4_x595),
.W_5(W_5_x595),
.W_6(W_6_x595),
.W_7(W_7_x595),
.W_8(W_8_x595),
.W_9(W_9_x595)
) u_28X28_x595 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x595),
 .score_0 (score_0_x595),
 .score_1 (score_1_x595),
 .score_2 (score_2_x595),
 .score_3 (score_3_x595),
 .score_4 (score_4_x595),
 .score_5 (score_5_x595),
 .score_6 (score_6_x595),
 .score_7 (score_7_x595),
 .score_8 (score_8_x595),
 .score_9 (score_9_x595)
);
 
myram_28X28 #(
.ID(596),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x596),
.W_1(W_1_x596),
.W_2(W_2_x596),
.W_3(W_3_x596),
.W_4(W_4_x596),
.W_5(W_5_x596),
.W_6(W_6_x596),
.W_7(W_7_x596),
.W_8(W_8_x596),
.W_9(W_9_x596)
) u_28X28_x596 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x596),
 .score_0 (score_0_x596),
 .score_1 (score_1_x596),
 .score_2 (score_2_x596),
 .score_3 (score_3_x596),
 .score_4 (score_4_x596),
 .score_5 (score_5_x596),
 .score_6 (score_6_x596),
 .score_7 (score_7_x596),
 .score_8 (score_8_x596),
 .score_9 (score_9_x596)
);
 
myram_28X28 #(
.ID(597),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x597),
.W_1(W_1_x597),
.W_2(W_2_x597),
.W_3(W_3_x597),
.W_4(W_4_x597),
.W_5(W_5_x597),
.W_6(W_6_x597),
.W_7(W_7_x597),
.W_8(W_8_x597),
.W_9(W_9_x597)
) u_28X28_x597 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x597),
 .score_0 (score_0_x597),
 .score_1 (score_1_x597),
 .score_2 (score_2_x597),
 .score_3 (score_3_x597),
 .score_4 (score_4_x597),
 .score_5 (score_5_x597),
 .score_6 (score_6_x597),
 .score_7 (score_7_x597),
 .score_8 (score_8_x597),
 .score_9 (score_9_x597)
);
 
myram_28X28 #(
.ID(598),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x598),
.W_1(W_1_x598),
.W_2(W_2_x598),
.W_3(W_3_x598),
.W_4(W_4_x598),
.W_5(W_5_x598),
.W_6(W_6_x598),
.W_7(W_7_x598),
.W_8(W_8_x598),
.W_9(W_9_x598)
) u_28X28_x598 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x598),
 .score_0 (score_0_x598),
 .score_1 (score_1_x598),
 .score_2 (score_2_x598),
 .score_3 (score_3_x598),
 .score_4 (score_4_x598),
 .score_5 (score_5_x598),
 .score_6 (score_6_x598),
 .score_7 (score_7_x598),
 .score_8 (score_8_x598),
 .score_9 (score_9_x598)
);
 
myram_28X28 #(
.ID(599),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x599),
.W_1(W_1_x599),
.W_2(W_2_x599),
.W_3(W_3_x599),
.W_4(W_4_x599),
.W_5(W_5_x599),
.W_6(W_6_x599),
.W_7(W_7_x599),
.W_8(W_8_x599),
.W_9(W_9_x599)
) u_28X28_x599 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x599),
 .score_0 (score_0_x599),
 .score_1 (score_1_x599),
 .score_2 (score_2_x599),
 .score_3 (score_3_x599),
 .score_4 (score_4_x599),
 .score_5 (score_5_x599),
 .score_6 (score_6_x599),
 .score_7 (score_7_x599),
 .score_8 (score_8_x599),
 .score_9 (score_9_x599)
);
 
myram_28X28 #(
.ID(600),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x600),
.W_1(W_1_x600),
.W_2(W_2_x600),
.W_3(W_3_x600),
.W_4(W_4_x600),
.W_5(W_5_x600),
.W_6(W_6_x600),
.W_7(W_7_x600),
.W_8(W_8_x600),
.W_9(W_9_x600)
) u_28X28_x600 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x600),
 .score_0 (score_0_x600),
 .score_1 (score_1_x600),
 .score_2 (score_2_x600),
 .score_3 (score_3_x600),
 .score_4 (score_4_x600),
 .score_5 (score_5_x600),
 .score_6 (score_6_x600),
 .score_7 (score_7_x600),
 .score_8 (score_8_x600),
 .score_9 (score_9_x600)
);
 
myram_28X28 #(
.ID(601),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x601),
.W_1(W_1_x601),
.W_2(W_2_x601),
.W_3(W_3_x601),
.W_4(W_4_x601),
.W_5(W_5_x601),
.W_6(W_6_x601),
.W_7(W_7_x601),
.W_8(W_8_x601),
.W_9(W_9_x601)
) u_28X28_x601 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x601),
 .score_0 (score_0_x601),
 .score_1 (score_1_x601),
 .score_2 (score_2_x601),
 .score_3 (score_3_x601),
 .score_4 (score_4_x601),
 .score_5 (score_5_x601),
 .score_6 (score_6_x601),
 .score_7 (score_7_x601),
 .score_8 (score_8_x601),
 .score_9 (score_9_x601)
);
 
myram_28X28 #(
.ID(602),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x602),
.W_1(W_1_x602),
.W_2(W_2_x602),
.W_3(W_3_x602),
.W_4(W_4_x602),
.W_5(W_5_x602),
.W_6(W_6_x602),
.W_7(W_7_x602),
.W_8(W_8_x602),
.W_9(W_9_x602)
) u_28X28_x602 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x602),
 .score_0 (score_0_x602),
 .score_1 (score_1_x602),
 .score_2 (score_2_x602),
 .score_3 (score_3_x602),
 .score_4 (score_4_x602),
 .score_5 (score_5_x602),
 .score_6 (score_6_x602),
 .score_7 (score_7_x602),
 .score_8 (score_8_x602),
 .score_9 (score_9_x602)
);
 
myram_28X28 #(
.ID(603),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x603),
.W_1(W_1_x603),
.W_2(W_2_x603),
.W_3(W_3_x603),
.W_4(W_4_x603),
.W_5(W_5_x603),
.W_6(W_6_x603),
.W_7(W_7_x603),
.W_8(W_8_x603),
.W_9(W_9_x603)
) u_28X28_x603 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x603),
 .score_0 (score_0_x603),
 .score_1 (score_1_x603),
 .score_2 (score_2_x603),
 .score_3 (score_3_x603),
 .score_4 (score_4_x603),
 .score_5 (score_5_x603),
 .score_6 (score_6_x603),
 .score_7 (score_7_x603),
 .score_8 (score_8_x603),
 .score_9 (score_9_x603)
);
 
myram_28X28 #(
.ID(604),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x604),
.W_1(W_1_x604),
.W_2(W_2_x604),
.W_3(W_3_x604),
.W_4(W_4_x604),
.W_5(W_5_x604),
.W_6(W_6_x604),
.W_7(W_7_x604),
.W_8(W_8_x604),
.W_9(W_9_x604)
) u_28X28_x604 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x604),
 .score_0 (score_0_x604),
 .score_1 (score_1_x604),
 .score_2 (score_2_x604),
 .score_3 (score_3_x604),
 .score_4 (score_4_x604),
 .score_5 (score_5_x604),
 .score_6 (score_6_x604),
 .score_7 (score_7_x604),
 .score_8 (score_8_x604),
 .score_9 (score_9_x604)
);
 
myram_28X28 #(
.ID(605),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x605),
.W_1(W_1_x605),
.W_2(W_2_x605),
.W_3(W_3_x605),
.W_4(W_4_x605),
.W_5(W_5_x605),
.W_6(W_6_x605),
.W_7(W_7_x605),
.W_8(W_8_x605),
.W_9(W_9_x605)
) u_28X28_x605 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x605),
 .score_0 (score_0_x605),
 .score_1 (score_1_x605),
 .score_2 (score_2_x605),
 .score_3 (score_3_x605),
 .score_4 (score_4_x605),
 .score_5 (score_5_x605),
 .score_6 (score_6_x605),
 .score_7 (score_7_x605),
 .score_8 (score_8_x605),
 .score_9 (score_9_x605)
);
 
myram_28X28 #(
.ID(606),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x606),
.W_1(W_1_x606),
.W_2(W_2_x606),
.W_3(W_3_x606),
.W_4(W_4_x606),
.W_5(W_5_x606),
.W_6(W_6_x606),
.W_7(W_7_x606),
.W_8(W_8_x606),
.W_9(W_9_x606)
) u_28X28_x606 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x606),
 .score_0 (score_0_x606),
 .score_1 (score_1_x606),
 .score_2 (score_2_x606),
 .score_3 (score_3_x606),
 .score_4 (score_4_x606),
 .score_5 (score_5_x606),
 .score_6 (score_6_x606),
 .score_7 (score_7_x606),
 .score_8 (score_8_x606),
 .score_9 (score_9_x606)
);
 
myram_28X28 #(
.ID(607),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x607),
.W_1(W_1_x607),
.W_2(W_2_x607),
.W_3(W_3_x607),
.W_4(W_4_x607),
.W_5(W_5_x607),
.W_6(W_6_x607),
.W_7(W_7_x607),
.W_8(W_8_x607),
.W_9(W_9_x607)
) u_28X28_x607 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x607),
 .score_0 (score_0_x607),
 .score_1 (score_1_x607),
 .score_2 (score_2_x607),
 .score_3 (score_3_x607),
 .score_4 (score_4_x607),
 .score_5 (score_5_x607),
 .score_6 (score_6_x607),
 .score_7 (score_7_x607),
 .score_8 (score_8_x607),
 .score_9 (score_9_x607)
);
 
myram_28X28 #(
.ID(608),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x608),
.W_1(W_1_x608),
.W_2(W_2_x608),
.W_3(W_3_x608),
.W_4(W_4_x608),
.W_5(W_5_x608),
.W_6(W_6_x608),
.W_7(W_7_x608),
.W_8(W_8_x608),
.W_9(W_9_x608)
) u_28X28_x608 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x608),
 .score_0 (score_0_x608),
 .score_1 (score_1_x608),
 .score_2 (score_2_x608),
 .score_3 (score_3_x608),
 .score_4 (score_4_x608),
 .score_5 (score_5_x608),
 .score_6 (score_6_x608),
 .score_7 (score_7_x608),
 .score_8 (score_8_x608),
 .score_9 (score_9_x608)
);
 
myram_28X28 #(
.ID(609),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x609),
.W_1(W_1_x609),
.W_2(W_2_x609),
.W_3(W_3_x609),
.W_4(W_4_x609),
.W_5(W_5_x609),
.W_6(W_6_x609),
.W_7(W_7_x609),
.W_8(W_8_x609),
.W_9(W_9_x609)
) u_28X28_x609 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x609),
 .score_0 (score_0_x609),
 .score_1 (score_1_x609),
 .score_2 (score_2_x609),
 .score_3 (score_3_x609),
 .score_4 (score_4_x609),
 .score_5 (score_5_x609),
 .score_6 (score_6_x609),
 .score_7 (score_7_x609),
 .score_8 (score_8_x609),
 .score_9 (score_9_x609)
);
 
myram_28X28 #(
.ID(610),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x610),
.W_1(W_1_x610),
.W_2(W_2_x610),
.W_3(W_3_x610),
.W_4(W_4_x610),
.W_5(W_5_x610),
.W_6(W_6_x610),
.W_7(W_7_x610),
.W_8(W_8_x610),
.W_9(W_9_x610)
) u_28X28_x610 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x610),
 .score_0 (score_0_x610),
 .score_1 (score_1_x610),
 .score_2 (score_2_x610),
 .score_3 (score_3_x610),
 .score_4 (score_4_x610),
 .score_5 (score_5_x610),
 .score_6 (score_6_x610),
 .score_7 (score_7_x610),
 .score_8 (score_8_x610),
 .score_9 (score_9_x610)
);
 
myram_28X28 #(
.ID(611),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x611),
.W_1(W_1_x611),
.W_2(W_2_x611),
.W_3(W_3_x611),
.W_4(W_4_x611),
.W_5(W_5_x611),
.W_6(W_6_x611),
.W_7(W_7_x611),
.W_8(W_8_x611),
.W_9(W_9_x611)
) u_28X28_x611 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x611),
 .score_0 (score_0_x611),
 .score_1 (score_1_x611),
 .score_2 (score_2_x611),
 .score_3 (score_3_x611),
 .score_4 (score_4_x611),
 .score_5 (score_5_x611),
 .score_6 (score_6_x611),
 .score_7 (score_7_x611),
 .score_8 (score_8_x611),
 .score_9 (score_9_x611)
);
 
myram_28X28 #(
.ID(612),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x612),
.W_1(W_1_x612),
.W_2(W_2_x612),
.W_3(W_3_x612),
.W_4(W_4_x612),
.W_5(W_5_x612),
.W_6(W_6_x612),
.W_7(W_7_x612),
.W_8(W_8_x612),
.W_9(W_9_x612)
) u_28X28_x612 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x612),
 .score_0 (score_0_x612),
 .score_1 (score_1_x612),
 .score_2 (score_2_x612),
 .score_3 (score_3_x612),
 .score_4 (score_4_x612),
 .score_5 (score_5_x612),
 .score_6 (score_6_x612),
 .score_7 (score_7_x612),
 .score_8 (score_8_x612),
 .score_9 (score_9_x612)
);
 
myram_28X28 #(
.ID(613),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x613),
.W_1(W_1_x613),
.W_2(W_2_x613),
.W_3(W_3_x613),
.W_4(W_4_x613),
.W_5(W_5_x613),
.W_6(W_6_x613),
.W_7(W_7_x613),
.W_8(W_8_x613),
.W_9(W_9_x613)
) u_28X28_x613 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x613),
 .score_0 (score_0_x613),
 .score_1 (score_1_x613),
 .score_2 (score_2_x613),
 .score_3 (score_3_x613),
 .score_4 (score_4_x613),
 .score_5 (score_5_x613),
 .score_6 (score_6_x613),
 .score_7 (score_7_x613),
 .score_8 (score_8_x613),
 .score_9 (score_9_x613)
);
 
myram_28X28 #(
.ID(614),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x614),
.W_1(W_1_x614),
.W_2(W_2_x614),
.W_3(W_3_x614),
.W_4(W_4_x614),
.W_5(W_5_x614),
.W_6(W_6_x614),
.W_7(W_7_x614),
.W_8(W_8_x614),
.W_9(W_9_x614)
) u_28X28_x614 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x614),
 .score_0 (score_0_x614),
 .score_1 (score_1_x614),
 .score_2 (score_2_x614),
 .score_3 (score_3_x614),
 .score_4 (score_4_x614),
 .score_5 (score_5_x614),
 .score_6 (score_6_x614),
 .score_7 (score_7_x614),
 .score_8 (score_8_x614),
 .score_9 (score_9_x614)
);
 
myram_28X28 #(
.ID(615),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x615),
.W_1(W_1_x615),
.W_2(W_2_x615),
.W_3(W_3_x615),
.W_4(W_4_x615),
.W_5(W_5_x615),
.W_6(W_6_x615),
.W_7(W_7_x615),
.W_8(W_8_x615),
.W_9(W_9_x615)
) u_28X28_x615 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x615),
 .score_0 (score_0_x615),
 .score_1 (score_1_x615),
 .score_2 (score_2_x615),
 .score_3 (score_3_x615),
 .score_4 (score_4_x615),
 .score_5 (score_5_x615),
 .score_6 (score_6_x615),
 .score_7 (score_7_x615),
 .score_8 (score_8_x615),
 .score_9 (score_9_x615)
);
 
myram_28X28 #(
.ID(616),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x616),
.W_1(W_1_x616),
.W_2(W_2_x616),
.W_3(W_3_x616),
.W_4(W_4_x616),
.W_5(W_5_x616),
.W_6(W_6_x616),
.W_7(W_7_x616),
.W_8(W_8_x616),
.W_9(W_9_x616)
) u_28X28_x616 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x616),
 .score_0 (score_0_x616),
 .score_1 (score_1_x616),
 .score_2 (score_2_x616),
 .score_3 (score_3_x616),
 .score_4 (score_4_x616),
 .score_5 (score_5_x616),
 .score_6 (score_6_x616),
 .score_7 (score_7_x616),
 .score_8 (score_8_x616),
 .score_9 (score_9_x616)
);
 
myram_28X28 #(
.ID(617),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x617),
.W_1(W_1_x617),
.W_2(W_2_x617),
.W_3(W_3_x617),
.W_4(W_4_x617),
.W_5(W_5_x617),
.W_6(W_6_x617),
.W_7(W_7_x617),
.W_8(W_8_x617),
.W_9(W_9_x617)
) u_28X28_x617 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x617),
 .score_0 (score_0_x617),
 .score_1 (score_1_x617),
 .score_2 (score_2_x617),
 .score_3 (score_3_x617),
 .score_4 (score_4_x617),
 .score_5 (score_5_x617),
 .score_6 (score_6_x617),
 .score_7 (score_7_x617),
 .score_8 (score_8_x617),
 .score_9 (score_9_x617)
);
 
myram_28X28 #(
.ID(618),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x618),
.W_1(W_1_x618),
.W_2(W_2_x618),
.W_3(W_3_x618),
.W_4(W_4_x618),
.W_5(W_5_x618),
.W_6(W_6_x618),
.W_7(W_7_x618),
.W_8(W_8_x618),
.W_9(W_9_x618)
) u_28X28_x618 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x618),
 .score_0 (score_0_x618),
 .score_1 (score_1_x618),
 .score_2 (score_2_x618),
 .score_3 (score_3_x618),
 .score_4 (score_4_x618),
 .score_5 (score_5_x618),
 .score_6 (score_6_x618),
 .score_7 (score_7_x618),
 .score_8 (score_8_x618),
 .score_9 (score_9_x618)
);
 
myram_28X28 #(
.ID(619),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x619),
.W_1(W_1_x619),
.W_2(W_2_x619),
.W_3(W_3_x619),
.W_4(W_4_x619),
.W_5(W_5_x619),
.W_6(W_6_x619),
.W_7(W_7_x619),
.W_8(W_8_x619),
.W_9(W_9_x619)
) u_28X28_x619 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x619),
 .score_0 (score_0_x619),
 .score_1 (score_1_x619),
 .score_2 (score_2_x619),
 .score_3 (score_3_x619),
 .score_4 (score_4_x619),
 .score_5 (score_5_x619),
 .score_6 (score_6_x619),
 .score_7 (score_7_x619),
 .score_8 (score_8_x619),
 .score_9 (score_9_x619)
);
 
myram_28X28 #(
.ID(620),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x620),
.W_1(W_1_x620),
.W_2(W_2_x620),
.W_3(W_3_x620),
.W_4(W_4_x620),
.W_5(W_5_x620),
.W_6(W_6_x620),
.W_7(W_7_x620),
.W_8(W_8_x620),
.W_9(W_9_x620)
) u_28X28_x620 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x620),
 .score_0 (score_0_x620),
 .score_1 (score_1_x620),
 .score_2 (score_2_x620),
 .score_3 (score_3_x620),
 .score_4 (score_4_x620),
 .score_5 (score_5_x620),
 .score_6 (score_6_x620),
 .score_7 (score_7_x620),
 .score_8 (score_8_x620),
 .score_9 (score_9_x620)
);
 
myram_28X28 #(
.ID(621),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x621),
.W_1(W_1_x621),
.W_2(W_2_x621),
.W_3(W_3_x621),
.W_4(W_4_x621),
.W_5(W_5_x621),
.W_6(W_6_x621),
.W_7(W_7_x621),
.W_8(W_8_x621),
.W_9(W_9_x621)
) u_28X28_x621 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x621),
 .score_0 (score_0_x621),
 .score_1 (score_1_x621),
 .score_2 (score_2_x621),
 .score_3 (score_3_x621),
 .score_4 (score_4_x621),
 .score_5 (score_5_x621),
 .score_6 (score_6_x621),
 .score_7 (score_7_x621),
 .score_8 (score_8_x621),
 .score_9 (score_9_x621)
);
 
myram_28X28 #(
.ID(622),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x622),
.W_1(W_1_x622),
.W_2(W_2_x622),
.W_3(W_3_x622),
.W_4(W_4_x622),
.W_5(W_5_x622),
.W_6(W_6_x622),
.W_7(W_7_x622),
.W_8(W_8_x622),
.W_9(W_9_x622)
) u_28X28_x622 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x622),
 .score_0 (score_0_x622),
 .score_1 (score_1_x622),
 .score_2 (score_2_x622),
 .score_3 (score_3_x622),
 .score_4 (score_4_x622),
 .score_5 (score_5_x622),
 .score_6 (score_6_x622),
 .score_7 (score_7_x622),
 .score_8 (score_8_x622),
 .score_9 (score_9_x622)
);
 
myram_28X28 #(
.ID(623),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x623),
.W_1(W_1_x623),
.W_2(W_2_x623),
.W_3(W_3_x623),
.W_4(W_4_x623),
.W_5(W_5_x623),
.W_6(W_6_x623),
.W_7(W_7_x623),
.W_8(W_8_x623),
.W_9(W_9_x623)
) u_28X28_x623 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x623),
 .score_0 (score_0_x623),
 .score_1 (score_1_x623),
 .score_2 (score_2_x623),
 .score_3 (score_3_x623),
 .score_4 (score_4_x623),
 .score_5 (score_5_x623),
 .score_6 (score_6_x623),
 .score_7 (score_7_x623),
 .score_8 (score_8_x623),
 .score_9 (score_9_x623)
);
 
myram_28X28 #(
.ID(624),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x624),
.W_1(W_1_x624),
.W_2(W_2_x624),
.W_3(W_3_x624),
.W_4(W_4_x624),
.W_5(W_5_x624),
.W_6(W_6_x624),
.W_7(W_7_x624),
.W_8(W_8_x624),
.W_9(W_9_x624)
) u_28X28_x624 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x624),
 .score_0 (score_0_x624),
 .score_1 (score_1_x624),
 .score_2 (score_2_x624),
 .score_3 (score_3_x624),
 .score_4 (score_4_x624),
 .score_5 (score_5_x624),
 .score_6 (score_6_x624),
 .score_7 (score_7_x624),
 .score_8 (score_8_x624),
 .score_9 (score_9_x624)
);
 
myram_28X28 #(
.ID(625),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x625),
.W_1(W_1_x625),
.W_2(W_2_x625),
.W_3(W_3_x625),
.W_4(W_4_x625),
.W_5(W_5_x625),
.W_6(W_6_x625),
.W_7(W_7_x625),
.W_8(W_8_x625),
.W_9(W_9_x625)
) u_28X28_x625 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x625),
 .score_0 (score_0_x625),
 .score_1 (score_1_x625),
 .score_2 (score_2_x625),
 .score_3 (score_3_x625),
 .score_4 (score_4_x625),
 .score_5 (score_5_x625),
 .score_6 (score_6_x625),
 .score_7 (score_7_x625),
 .score_8 (score_8_x625),
 .score_9 (score_9_x625)
);
 
myram_28X28 #(
.ID(626),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x626),
.W_1(W_1_x626),
.W_2(W_2_x626),
.W_3(W_3_x626),
.W_4(W_4_x626),
.W_5(W_5_x626),
.W_6(W_6_x626),
.W_7(W_7_x626),
.W_8(W_8_x626),
.W_9(W_9_x626)
) u_28X28_x626 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x626),
 .score_0 (score_0_x626),
 .score_1 (score_1_x626),
 .score_2 (score_2_x626),
 .score_3 (score_3_x626),
 .score_4 (score_4_x626),
 .score_5 (score_5_x626),
 .score_6 (score_6_x626),
 .score_7 (score_7_x626),
 .score_8 (score_8_x626),
 .score_9 (score_9_x626)
);
 
myram_28X28 #(
.ID(627),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x627),
.W_1(W_1_x627),
.W_2(W_2_x627),
.W_3(W_3_x627),
.W_4(W_4_x627),
.W_5(W_5_x627),
.W_6(W_6_x627),
.W_7(W_7_x627),
.W_8(W_8_x627),
.W_9(W_9_x627)
) u_28X28_x627 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x627),
 .score_0 (score_0_x627),
 .score_1 (score_1_x627),
 .score_2 (score_2_x627),
 .score_3 (score_3_x627),
 .score_4 (score_4_x627),
 .score_5 (score_5_x627),
 .score_6 (score_6_x627),
 .score_7 (score_7_x627),
 .score_8 (score_8_x627),
 .score_9 (score_9_x627)
);
 
myram_28X28 #(
.ID(628),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x628),
.W_1(W_1_x628),
.W_2(W_2_x628),
.W_3(W_3_x628),
.W_4(W_4_x628),
.W_5(W_5_x628),
.W_6(W_6_x628),
.W_7(W_7_x628),
.W_8(W_8_x628),
.W_9(W_9_x628)
) u_28X28_x628 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x628),
 .score_0 (score_0_x628),
 .score_1 (score_1_x628),
 .score_2 (score_2_x628),
 .score_3 (score_3_x628),
 .score_4 (score_4_x628),
 .score_5 (score_5_x628),
 .score_6 (score_6_x628),
 .score_7 (score_7_x628),
 .score_8 (score_8_x628),
 .score_9 (score_9_x628)
);
 
myram_28X28 #(
.ID(629),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x629),
.W_1(W_1_x629),
.W_2(W_2_x629),
.W_3(W_3_x629),
.W_4(W_4_x629),
.W_5(W_5_x629),
.W_6(W_6_x629),
.W_7(W_7_x629),
.W_8(W_8_x629),
.W_9(W_9_x629)
) u_28X28_x629 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x629),
 .score_0 (score_0_x629),
 .score_1 (score_1_x629),
 .score_2 (score_2_x629),
 .score_3 (score_3_x629),
 .score_4 (score_4_x629),
 .score_5 (score_5_x629),
 .score_6 (score_6_x629),
 .score_7 (score_7_x629),
 .score_8 (score_8_x629),
 .score_9 (score_9_x629)
);
 
myram_28X28 #(
.ID(630),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x630),
.W_1(W_1_x630),
.W_2(W_2_x630),
.W_3(W_3_x630),
.W_4(W_4_x630),
.W_5(W_5_x630),
.W_6(W_6_x630),
.W_7(W_7_x630),
.W_8(W_8_x630),
.W_9(W_9_x630)
) u_28X28_x630 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x630),
 .score_0 (score_0_x630),
 .score_1 (score_1_x630),
 .score_2 (score_2_x630),
 .score_3 (score_3_x630),
 .score_4 (score_4_x630),
 .score_5 (score_5_x630),
 .score_6 (score_6_x630),
 .score_7 (score_7_x630),
 .score_8 (score_8_x630),
 .score_9 (score_9_x630)
);
 
myram_28X28 #(
.ID(631),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x631),
.W_1(W_1_x631),
.W_2(W_2_x631),
.W_3(W_3_x631),
.W_4(W_4_x631),
.W_5(W_5_x631),
.W_6(W_6_x631),
.W_7(W_7_x631),
.W_8(W_8_x631),
.W_9(W_9_x631)
) u_28X28_x631 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x631),
 .score_0 (score_0_x631),
 .score_1 (score_1_x631),
 .score_2 (score_2_x631),
 .score_3 (score_3_x631),
 .score_4 (score_4_x631),
 .score_5 (score_5_x631),
 .score_6 (score_6_x631),
 .score_7 (score_7_x631),
 .score_8 (score_8_x631),
 .score_9 (score_9_x631)
);
 
myram_28X28 #(
.ID(632),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x632),
.W_1(W_1_x632),
.W_2(W_2_x632),
.W_3(W_3_x632),
.W_4(W_4_x632),
.W_5(W_5_x632),
.W_6(W_6_x632),
.W_7(W_7_x632),
.W_8(W_8_x632),
.W_9(W_9_x632)
) u_28X28_x632 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x632),
 .score_0 (score_0_x632),
 .score_1 (score_1_x632),
 .score_2 (score_2_x632),
 .score_3 (score_3_x632),
 .score_4 (score_4_x632),
 .score_5 (score_5_x632),
 .score_6 (score_6_x632),
 .score_7 (score_7_x632),
 .score_8 (score_8_x632),
 .score_9 (score_9_x632)
);
 
myram_28X28 #(
.ID(633),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x633),
.W_1(W_1_x633),
.W_2(W_2_x633),
.W_3(W_3_x633),
.W_4(W_4_x633),
.W_5(W_5_x633),
.W_6(W_6_x633),
.W_7(W_7_x633),
.W_8(W_8_x633),
.W_9(W_9_x633)
) u_28X28_x633 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x633),
 .score_0 (score_0_x633),
 .score_1 (score_1_x633),
 .score_2 (score_2_x633),
 .score_3 (score_3_x633),
 .score_4 (score_4_x633),
 .score_5 (score_5_x633),
 .score_6 (score_6_x633),
 .score_7 (score_7_x633),
 .score_8 (score_8_x633),
 .score_9 (score_9_x633)
);
 
myram_28X28 #(
.ID(634),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x634),
.W_1(W_1_x634),
.W_2(W_2_x634),
.W_3(W_3_x634),
.W_4(W_4_x634),
.W_5(W_5_x634),
.W_6(W_6_x634),
.W_7(W_7_x634),
.W_8(W_8_x634),
.W_9(W_9_x634)
) u_28X28_x634 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x634),
 .score_0 (score_0_x634),
 .score_1 (score_1_x634),
 .score_2 (score_2_x634),
 .score_3 (score_3_x634),
 .score_4 (score_4_x634),
 .score_5 (score_5_x634),
 .score_6 (score_6_x634),
 .score_7 (score_7_x634),
 .score_8 (score_8_x634),
 .score_9 (score_9_x634)
);
 
myram_28X28 #(
.ID(635),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x635),
.W_1(W_1_x635),
.W_2(W_2_x635),
.W_3(W_3_x635),
.W_4(W_4_x635),
.W_5(W_5_x635),
.W_6(W_6_x635),
.W_7(W_7_x635),
.W_8(W_8_x635),
.W_9(W_9_x635)
) u_28X28_x635 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x635),
 .score_0 (score_0_x635),
 .score_1 (score_1_x635),
 .score_2 (score_2_x635),
 .score_3 (score_3_x635),
 .score_4 (score_4_x635),
 .score_5 (score_5_x635),
 .score_6 (score_6_x635),
 .score_7 (score_7_x635),
 .score_8 (score_8_x635),
 .score_9 (score_9_x635)
);
 
myram_28X28 #(
.ID(636),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x636),
.W_1(W_1_x636),
.W_2(W_2_x636),
.W_3(W_3_x636),
.W_4(W_4_x636),
.W_5(W_5_x636),
.W_6(W_6_x636),
.W_7(W_7_x636),
.W_8(W_8_x636),
.W_9(W_9_x636)
) u_28X28_x636 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x636),
 .score_0 (score_0_x636),
 .score_1 (score_1_x636),
 .score_2 (score_2_x636),
 .score_3 (score_3_x636),
 .score_4 (score_4_x636),
 .score_5 (score_5_x636),
 .score_6 (score_6_x636),
 .score_7 (score_7_x636),
 .score_8 (score_8_x636),
 .score_9 (score_9_x636)
);
 
myram_28X28 #(
.ID(637),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x637),
.W_1(W_1_x637),
.W_2(W_2_x637),
.W_3(W_3_x637),
.W_4(W_4_x637),
.W_5(W_5_x637),
.W_6(W_6_x637),
.W_7(W_7_x637),
.W_8(W_8_x637),
.W_9(W_9_x637)
) u_28X28_x637 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x637),
 .score_0 (score_0_x637),
 .score_1 (score_1_x637),
 .score_2 (score_2_x637),
 .score_3 (score_3_x637),
 .score_4 (score_4_x637),
 .score_5 (score_5_x637),
 .score_6 (score_6_x637),
 .score_7 (score_7_x637),
 .score_8 (score_8_x637),
 .score_9 (score_9_x637)
);
 
myram_28X28 #(
.ID(638),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x638),
.W_1(W_1_x638),
.W_2(W_2_x638),
.W_3(W_3_x638),
.W_4(W_4_x638),
.W_5(W_5_x638),
.W_6(W_6_x638),
.W_7(W_7_x638),
.W_8(W_8_x638),
.W_9(W_9_x638)
) u_28X28_x638 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x638),
 .score_0 (score_0_x638),
 .score_1 (score_1_x638),
 .score_2 (score_2_x638),
 .score_3 (score_3_x638),
 .score_4 (score_4_x638),
 .score_5 (score_5_x638),
 .score_6 (score_6_x638),
 .score_7 (score_7_x638),
 .score_8 (score_8_x638),
 .score_9 (score_9_x638)
);
 
myram_28X28 #(
.ID(639),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x639),
.W_1(W_1_x639),
.W_2(W_2_x639),
.W_3(W_3_x639),
.W_4(W_4_x639),
.W_5(W_5_x639),
.W_6(W_6_x639),
.W_7(W_7_x639),
.W_8(W_8_x639),
.W_9(W_9_x639)
) u_28X28_x639 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x639),
 .score_0 (score_0_x639),
 .score_1 (score_1_x639),
 .score_2 (score_2_x639),
 .score_3 (score_3_x639),
 .score_4 (score_4_x639),
 .score_5 (score_5_x639),
 .score_6 (score_6_x639),
 .score_7 (score_7_x639),
 .score_8 (score_8_x639),
 .score_9 (score_9_x639)
);
 
myram_28X28 #(
.ID(640),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x640),
.W_1(W_1_x640),
.W_2(W_2_x640),
.W_3(W_3_x640),
.W_4(W_4_x640),
.W_5(W_5_x640),
.W_6(W_6_x640),
.W_7(W_7_x640),
.W_8(W_8_x640),
.W_9(W_9_x640)
) u_28X28_x640 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x640),
 .score_0 (score_0_x640),
 .score_1 (score_1_x640),
 .score_2 (score_2_x640),
 .score_3 (score_3_x640),
 .score_4 (score_4_x640),
 .score_5 (score_5_x640),
 .score_6 (score_6_x640),
 .score_7 (score_7_x640),
 .score_8 (score_8_x640),
 .score_9 (score_9_x640)
);
 
myram_28X28 #(
.ID(641),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x641),
.W_1(W_1_x641),
.W_2(W_2_x641),
.W_3(W_3_x641),
.W_4(W_4_x641),
.W_5(W_5_x641),
.W_6(W_6_x641),
.W_7(W_7_x641),
.W_8(W_8_x641),
.W_9(W_9_x641)
) u_28X28_x641 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x641),
 .score_0 (score_0_x641),
 .score_1 (score_1_x641),
 .score_2 (score_2_x641),
 .score_3 (score_3_x641),
 .score_4 (score_4_x641),
 .score_5 (score_5_x641),
 .score_6 (score_6_x641),
 .score_7 (score_7_x641),
 .score_8 (score_8_x641),
 .score_9 (score_9_x641)
);
 
myram_28X28 #(
.ID(642),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x642),
.W_1(W_1_x642),
.W_2(W_2_x642),
.W_3(W_3_x642),
.W_4(W_4_x642),
.W_5(W_5_x642),
.W_6(W_6_x642),
.W_7(W_7_x642),
.W_8(W_8_x642),
.W_9(W_9_x642)
) u_28X28_x642 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x642),
 .score_0 (score_0_x642),
 .score_1 (score_1_x642),
 .score_2 (score_2_x642),
 .score_3 (score_3_x642),
 .score_4 (score_4_x642),
 .score_5 (score_5_x642),
 .score_6 (score_6_x642),
 .score_7 (score_7_x642),
 .score_8 (score_8_x642),
 .score_9 (score_9_x642)
);
 
myram_28X28 #(
.ID(643),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x643),
.W_1(W_1_x643),
.W_2(W_2_x643),
.W_3(W_3_x643),
.W_4(W_4_x643),
.W_5(W_5_x643),
.W_6(W_6_x643),
.W_7(W_7_x643),
.W_8(W_8_x643),
.W_9(W_9_x643)
) u_28X28_x643 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x643),
 .score_0 (score_0_x643),
 .score_1 (score_1_x643),
 .score_2 (score_2_x643),
 .score_3 (score_3_x643),
 .score_4 (score_4_x643),
 .score_5 (score_5_x643),
 .score_6 (score_6_x643),
 .score_7 (score_7_x643),
 .score_8 (score_8_x643),
 .score_9 (score_9_x643)
);
 
myram_28X28 #(
.ID(644),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x644),
.W_1(W_1_x644),
.W_2(W_2_x644),
.W_3(W_3_x644),
.W_4(W_4_x644),
.W_5(W_5_x644),
.W_6(W_6_x644),
.W_7(W_7_x644),
.W_8(W_8_x644),
.W_9(W_9_x644)
) u_28X28_x644 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x644),
 .score_0 (score_0_x644),
 .score_1 (score_1_x644),
 .score_2 (score_2_x644),
 .score_3 (score_3_x644),
 .score_4 (score_4_x644),
 .score_5 (score_5_x644),
 .score_6 (score_6_x644),
 .score_7 (score_7_x644),
 .score_8 (score_8_x644),
 .score_9 (score_9_x644)
);
 
myram_28X28 #(
.ID(645),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x645),
.W_1(W_1_x645),
.W_2(W_2_x645),
.W_3(W_3_x645),
.W_4(W_4_x645),
.W_5(W_5_x645),
.W_6(W_6_x645),
.W_7(W_7_x645),
.W_8(W_8_x645),
.W_9(W_9_x645)
) u_28X28_x645 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x645),
 .score_0 (score_0_x645),
 .score_1 (score_1_x645),
 .score_2 (score_2_x645),
 .score_3 (score_3_x645),
 .score_4 (score_4_x645),
 .score_5 (score_5_x645),
 .score_6 (score_6_x645),
 .score_7 (score_7_x645),
 .score_8 (score_8_x645),
 .score_9 (score_9_x645)
);
 
myram_28X28 #(
.ID(646),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x646),
.W_1(W_1_x646),
.W_2(W_2_x646),
.W_3(W_3_x646),
.W_4(W_4_x646),
.W_5(W_5_x646),
.W_6(W_6_x646),
.W_7(W_7_x646),
.W_8(W_8_x646),
.W_9(W_9_x646)
) u_28X28_x646 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x646),
 .score_0 (score_0_x646),
 .score_1 (score_1_x646),
 .score_2 (score_2_x646),
 .score_3 (score_3_x646),
 .score_4 (score_4_x646),
 .score_5 (score_5_x646),
 .score_6 (score_6_x646),
 .score_7 (score_7_x646),
 .score_8 (score_8_x646),
 .score_9 (score_9_x646)
);
 
myram_28X28 #(
.ID(647),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x647),
.W_1(W_1_x647),
.W_2(W_2_x647),
.W_3(W_3_x647),
.W_4(W_4_x647),
.W_5(W_5_x647),
.W_6(W_6_x647),
.W_7(W_7_x647),
.W_8(W_8_x647),
.W_9(W_9_x647)
) u_28X28_x647 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x647),
 .score_0 (score_0_x647),
 .score_1 (score_1_x647),
 .score_2 (score_2_x647),
 .score_3 (score_3_x647),
 .score_4 (score_4_x647),
 .score_5 (score_5_x647),
 .score_6 (score_6_x647),
 .score_7 (score_7_x647),
 .score_8 (score_8_x647),
 .score_9 (score_9_x647)
);
 
myram_28X28 #(
.ID(648),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x648),
.W_1(W_1_x648),
.W_2(W_2_x648),
.W_3(W_3_x648),
.W_4(W_4_x648),
.W_5(W_5_x648),
.W_6(W_6_x648),
.W_7(W_7_x648),
.W_8(W_8_x648),
.W_9(W_9_x648)
) u_28X28_x648 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x648),
 .score_0 (score_0_x648),
 .score_1 (score_1_x648),
 .score_2 (score_2_x648),
 .score_3 (score_3_x648),
 .score_4 (score_4_x648),
 .score_5 (score_5_x648),
 .score_6 (score_6_x648),
 .score_7 (score_7_x648),
 .score_8 (score_8_x648),
 .score_9 (score_9_x648)
);
 
myram_28X28 #(
.ID(649),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x649),
.W_1(W_1_x649),
.W_2(W_2_x649),
.W_3(W_3_x649),
.W_4(W_4_x649),
.W_5(W_5_x649),
.W_6(W_6_x649),
.W_7(W_7_x649),
.W_8(W_8_x649),
.W_9(W_9_x649)
) u_28X28_x649 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x649),
 .score_0 (score_0_x649),
 .score_1 (score_1_x649),
 .score_2 (score_2_x649),
 .score_3 (score_3_x649),
 .score_4 (score_4_x649),
 .score_5 (score_5_x649),
 .score_6 (score_6_x649),
 .score_7 (score_7_x649),
 .score_8 (score_8_x649),
 .score_9 (score_9_x649)
);
 
myram_28X28 #(
.ID(650),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x650),
.W_1(W_1_x650),
.W_2(W_2_x650),
.W_3(W_3_x650),
.W_4(W_4_x650),
.W_5(W_5_x650),
.W_6(W_6_x650),
.W_7(W_7_x650),
.W_8(W_8_x650),
.W_9(W_9_x650)
) u_28X28_x650 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x650),
 .score_0 (score_0_x650),
 .score_1 (score_1_x650),
 .score_2 (score_2_x650),
 .score_3 (score_3_x650),
 .score_4 (score_4_x650),
 .score_5 (score_5_x650),
 .score_6 (score_6_x650),
 .score_7 (score_7_x650),
 .score_8 (score_8_x650),
 .score_9 (score_9_x650)
);
 
myram_28X28 #(
.ID(651),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x651),
.W_1(W_1_x651),
.W_2(W_2_x651),
.W_3(W_3_x651),
.W_4(W_4_x651),
.W_5(W_5_x651),
.W_6(W_6_x651),
.W_7(W_7_x651),
.W_8(W_8_x651),
.W_9(W_9_x651)
) u_28X28_x651 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x651),
 .score_0 (score_0_x651),
 .score_1 (score_1_x651),
 .score_2 (score_2_x651),
 .score_3 (score_3_x651),
 .score_4 (score_4_x651),
 .score_5 (score_5_x651),
 .score_6 (score_6_x651),
 .score_7 (score_7_x651),
 .score_8 (score_8_x651),
 .score_9 (score_9_x651)
);
 
myram_28X28 #(
.ID(652),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x652),
.W_1(W_1_x652),
.W_2(W_2_x652),
.W_3(W_3_x652),
.W_4(W_4_x652),
.W_5(W_5_x652),
.W_6(W_6_x652),
.W_7(W_7_x652),
.W_8(W_8_x652),
.W_9(W_9_x652)
) u_28X28_x652 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x652),
 .score_0 (score_0_x652),
 .score_1 (score_1_x652),
 .score_2 (score_2_x652),
 .score_3 (score_3_x652),
 .score_4 (score_4_x652),
 .score_5 (score_5_x652),
 .score_6 (score_6_x652),
 .score_7 (score_7_x652),
 .score_8 (score_8_x652),
 .score_9 (score_9_x652)
);
 
myram_28X28 #(
.ID(653),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x653),
.W_1(W_1_x653),
.W_2(W_2_x653),
.W_3(W_3_x653),
.W_4(W_4_x653),
.W_5(W_5_x653),
.W_6(W_6_x653),
.W_7(W_7_x653),
.W_8(W_8_x653),
.W_9(W_9_x653)
) u_28X28_x653 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x653),
 .score_0 (score_0_x653),
 .score_1 (score_1_x653),
 .score_2 (score_2_x653),
 .score_3 (score_3_x653),
 .score_4 (score_4_x653),
 .score_5 (score_5_x653),
 .score_6 (score_6_x653),
 .score_7 (score_7_x653),
 .score_8 (score_8_x653),
 .score_9 (score_9_x653)
);
 
myram_28X28 #(
.ID(654),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x654),
.W_1(W_1_x654),
.W_2(W_2_x654),
.W_3(W_3_x654),
.W_4(W_4_x654),
.W_5(W_5_x654),
.W_6(W_6_x654),
.W_7(W_7_x654),
.W_8(W_8_x654),
.W_9(W_9_x654)
) u_28X28_x654 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x654),
 .score_0 (score_0_x654),
 .score_1 (score_1_x654),
 .score_2 (score_2_x654),
 .score_3 (score_3_x654),
 .score_4 (score_4_x654),
 .score_5 (score_5_x654),
 .score_6 (score_6_x654),
 .score_7 (score_7_x654),
 .score_8 (score_8_x654),
 .score_9 (score_9_x654)
);
 
myram_28X28 #(
.ID(655),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x655),
.W_1(W_1_x655),
.W_2(W_2_x655),
.W_3(W_3_x655),
.W_4(W_4_x655),
.W_5(W_5_x655),
.W_6(W_6_x655),
.W_7(W_7_x655),
.W_8(W_8_x655),
.W_9(W_9_x655)
) u_28X28_x655 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x655),
 .score_0 (score_0_x655),
 .score_1 (score_1_x655),
 .score_2 (score_2_x655),
 .score_3 (score_3_x655),
 .score_4 (score_4_x655),
 .score_5 (score_5_x655),
 .score_6 (score_6_x655),
 .score_7 (score_7_x655),
 .score_8 (score_8_x655),
 .score_9 (score_9_x655)
);
 
myram_28X28 #(
.ID(656),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x656),
.W_1(W_1_x656),
.W_2(W_2_x656),
.W_3(W_3_x656),
.W_4(W_4_x656),
.W_5(W_5_x656),
.W_6(W_6_x656),
.W_7(W_7_x656),
.W_8(W_8_x656),
.W_9(W_9_x656)
) u_28X28_x656 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x656),
 .score_0 (score_0_x656),
 .score_1 (score_1_x656),
 .score_2 (score_2_x656),
 .score_3 (score_3_x656),
 .score_4 (score_4_x656),
 .score_5 (score_5_x656),
 .score_6 (score_6_x656),
 .score_7 (score_7_x656),
 .score_8 (score_8_x656),
 .score_9 (score_9_x656)
);
 
myram_28X28 #(
.ID(657),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x657),
.W_1(W_1_x657),
.W_2(W_2_x657),
.W_3(W_3_x657),
.W_4(W_4_x657),
.W_5(W_5_x657),
.W_6(W_6_x657),
.W_7(W_7_x657),
.W_8(W_8_x657),
.W_9(W_9_x657)
) u_28X28_x657 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x657),
 .score_0 (score_0_x657),
 .score_1 (score_1_x657),
 .score_2 (score_2_x657),
 .score_3 (score_3_x657),
 .score_4 (score_4_x657),
 .score_5 (score_5_x657),
 .score_6 (score_6_x657),
 .score_7 (score_7_x657),
 .score_8 (score_8_x657),
 .score_9 (score_9_x657)
);
 
myram_28X28 #(
.ID(658),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x658),
.W_1(W_1_x658),
.W_2(W_2_x658),
.W_3(W_3_x658),
.W_4(W_4_x658),
.W_5(W_5_x658),
.W_6(W_6_x658),
.W_7(W_7_x658),
.W_8(W_8_x658),
.W_9(W_9_x658)
) u_28X28_x658 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x658),
 .score_0 (score_0_x658),
 .score_1 (score_1_x658),
 .score_2 (score_2_x658),
 .score_3 (score_3_x658),
 .score_4 (score_4_x658),
 .score_5 (score_5_x658),
 .score_6 (score_6_x658),
 .score_7 (score_7_x658),
 .score_8 (score_8_x658),
 .score_9 (score_9_x658)
);
 
myram_28X28 #(
.ID(659),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x659),
.W_1(W_1_x659),
.W_2(W_2_x659),
.W_3(W_3_x659),
.W_4(W_4_x659),
.W_5(W_5_x659),
.W_6(W_6_x659),
.W_7(W_7_x659),
.W_8(W_8_x659),
.W_9(W_9_x659)
) u_28X28_x659 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x659),
 .score_0 (score_0_x659),
 .score_1 (score_1_x659),
 .score_2 (score_2_x659),
 .score_3 (score_3_x659),
 .score_4 (score_4_x659),
 .score_5 (score_5_x659),
 .score_6 (score_6_x659),
 .score_7 (score_7_x659),
 .score_8 (score_8_x659),
 .score_9 (score_9_x659)
);
 
myram_28X28 #(
.ID(660),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x660),
.W_1(W_1_x660),
.W_2(W_2_x660),
.W_3(W_3_x660),
.W_4(W_4_x660),
.W_5(W_5_x660),
.W_6(W_6_x660),
.W_7(W_7_x660),
.W_8(W_8_x660),
.W_9(W_9_x660)
) u_28X28_x660 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x660),
 .score_0 (score_0_x660),
 .score_1 (score_1_x660),
 .score_2 (score_2_x660),
 .score_3 (score_3_x660),
 .score_4 (score_4_x660),
 .score_5 (score_5_x660),
 .score_6 (score_6_x660),
 .score_7 (score_7_x660),
 .score_8 (score_8_x660),
 .score_9 (score_9_x660)
);
 
myram_28X28 #(
.ID(661),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x661),
.W_1(W_1_x661),
.W_2(W_2_x661),
.W_3(W_3_x661),
.W_4(W_4_x661),
.W_5(W_5_x661),
.W_6(W_6_x661),
.W_7(W_7_x661),
.W_8(W_8_x661),
.W_9(W_9_x661)
) u_28X28_x661 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x661),
 .score_0 (score_0_x661),
 .score_1 (score_1_x661),
 .score_2 (score_2_x661),
 .score_3 (score_3_x661),
 .score_4 (score_4_x661),
 .score_5 (score_5_x661),
 .score_6 (score_6_x661),
 .score_7 (score_7_x661),
 .score_8 (score_8_x661),
 .score_9 (score_9_x661)
);
 
myram_28X28 #(
.ID(662),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x662),
.W_1(W_1_x662),
.W_2(W_2_x662),
.W_3(W_3_x662),
.W_4(W_4_x662),
.W_5(W_5_x662),
.W_6(W_6_x662),
.W_7(W_7_x662),
.W_8(W_8_x662),
.W_9(W_9_x662)
) u_28X28_x662 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x662),
 .score_0 (score_0_x662),
 .score_1 (score_1_x662),
 .score_2 (score_2_x662),
 .score_3 (score_3_x662),
 .score_4 (score_4_x662),
 .score_5 (score_5_x662),
 .score_6 (score_6_x662),
 .score_7 (score_7_x662),
 .score_8 (score_8_x662),
 .score_9 (score_9_x662)
);
 
myram_28X28 #(
.ID(663),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x663),
.W_1(W_1_x663),
.W_2(W_2_x663),
.W_3(W_3_x663),
.W_4(W_4_x663),
.W_5(W_5_x663),
.W_6(W_6_x663),
.W_7(W_7_x663),
.W_8(W_8_x663),
.W_9(W_9_x663)
) u_28X28_x663 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x663),
 .score_0 (score_0_x663),
 .score_1 (score_1_x663),
 .score_2 (score_2_x663),
 .score_3 (score_3_x663),
 .score_4 (score_4_x663),
 .score_5 (score_5_x663),
 .score_6 (score_6_x663),
 .score_7 (score_7_x663),
 .score_8 (score_8_x663),
 .score_9 (score_9_x663)
);
 
myram_28X28 #(
.ID(664),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x664),
.W_1(W_1_x664),
.W_2(W_2_x664),
.W_3(W_3_x664),
.W_4(W_4_x664),
.W_5(W_5_x664),
.W_6(W_6_x664),
.W_7(W_7_x664),
.W_8(W_8_x664),
.W_9(W_9_x664)
) u_28X28_x664 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x664),
 .score_0 (score_0_x664),
 .score_1 (score_1_x664),
 .score_2 (score_2_x664),
 .score_3 (score_3_x664),
 .score_4 (score_4_x664),
 .score_5 (score_5_x664),
 .score_6 (score_6_x664),
 .score_7 (score_7_x664),
 .score_8 (score_8_x664),
 .score_9 (score_9_x664)
);
 
myram_28X28 #(
.ID(665),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x665),
.W_1(W_1_x665),
.W_2(W_2_x665),
.W_3(W_3_x665),
.W_4(W_4_x665),
.W_5(W_5_x665),
.W_6(W_6_x665),
.W_7(W_7_x665),
.W_8(W_8_x665),
.W_9(W_9_x665)
) u_28X28_x665 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x665),
 .score_0 (score_0_x665),
 .score_1 (score_1_x665),
 .score_2 (score_2_x665),
 .score_3 (score_3_x665),
 .score_4 (score_4_x665),
 .score_5 (score_5_x665),
 .score_6 (score_6_x665),
 .score_7 (score_7_x665),
 .score_8 (score_8_x665),
 .score_9 (score_9_x665)
);
 
myram_28X28 #(
.ID(666),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x666),
.W_1(W_1_x666),
.W_2(W_2_x666),
.W_3(W_3_x666),
.W_4(W_4_x666),
.W_5(W_5_x666),
.W_6(W_6_x666),
.W_7(W_7_x666),
.W_8(W_8_x666),
.W_9(W_9_x666)
) u_28X28_x666 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x666),
 .score_0 (score_0_x666),
 .score_1 (score_1_x666),
 .score_2 (score_2_x666),
 .score_3 (score_3_x666),
 .score_4 (score_4_x666),
 .score_5 (score_5_x666),
 .score_6 (score_6_x666),
 .score_7 (score_7_x666),
 .score_8 (score_8_x666),
 .score_9 (score_9_x666)
);
 
myram_28X28 #(
.ID(667),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x667),
.W_1(W_1_x667),
.W_2(W_2_x667),
.W_3(W_3_x667),
.W_4(W_4_x667),
.W_5(W_5_x667),
.W_6(W_6_x667),
.W_7(W_7_x667),
.W_8(W_8_x667),
.W_9(W_9_x667)
) u_28X28_x667 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x667),
 .score_0 (score_0_x667),
 .score_1 (score_1_x667),
 .score_2 (score_2_x667),
 .score_3 (score_3_x667),
 .score_4 (score_4_x667),
 .score_5 (score_5_x667),
 .score_6 (score_6_x667),
 .score_7 (score_7_x667),
 .score_8 (score_8_x667),
 .score_9 (score_9_x667)
);
 
myram_28X28 #(
.ID(668),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x668),
.W_1(W_1_x668),
.W_2(W_2_x668),
.W_3(W_3_x668),
.W_4(W_4_x668),
.W_5(W_5_x668),
.W_6(W_6_x668),
.W_7(W_7_x668),
.W_8(W_8_x668),
.W_9(W_9_x668)
) u_28X28_x668 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x668),
 .score_0 (score_0_x668),
 .score_1 (score_1_x668),
 .score_2 (score_2_x668),
 .score_3 (score_3_x668),
 .score_4 (score_4_x668),
 .score_5 (score_5_x668),
 .score_6 (score_6_x668),
 .score_7 (score_7_x668),
 .score_8 (score_8_x668),
 .score_9 (score_9_x668)
);
 
myram_28X28 #(
.ID(669),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x669),
.W_1(W_1_x669),
.W_2(W_2_x669),
.W_3(W_3_x669),
.W_4(W_4_x669),
.W_5(W_5_x669),
.W_6(W_6_x669),
.W_7(W_7_x669),
.W_8(W_8_x669),
.W_9(W_9_x669)
) u_28X28_x669 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x669),
 .score_0 (score_0_x669),
 .score_1 (score_1_x669),
 .score_2 (score_2_x669),
 .score_3 (score_3_x669),
 .score_4 (score_4_x669),
 .score_5 (score_5_x669),
 .score_6 (score_6_x669),
 .score_7 (score_7_x669),
 .score_8 (score_8_x669),
 .score_9 (score_9_x669)
);
 
myram_28X28 #(
.ID(670),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x670),
.W_1(W_1_x670),
.W_2(W_2_x670),
.W_3(W_3_x670),
.W_4(W_4_x670),
.W_5(W_5_x670),
.W_6(W_6_x670),
.W_7(W_7_x670),
.W_8(W_8_x670),
.W_9(W_9_x670)
) u_28X28_x670 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x670),
 .score_0 (score_0_x670),
 .score_1 (score_1_x670),
 .score_2 (score_2_x670),
 .score_3 (score_3_x670),
 .score_4 (score_4_x670),
 .score_5 (score_5_x670),
 .score_6 (score_6_x670),
 .score_7 (score_7_x670),
 .score_8 (score_8_x670),
 .score_9 (score_9_x670)
);
 
myram_28X28 #(
.ID(671),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x671),
.W_1(W_1_x671),
.W_2(W_2_x671),
.W_3(W_3_x671),
.W_4(W_4_x671),
.W_5(W_5_x671),
.W_6(W_6_x671),
.W_7(W_7_x671),
.W_8(W_8_x671),
.W_9(W_9_x671)
) u_28X28_x671 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x671),
 .score_0 (score_0_x671),
 .score_1 (score_1_x671),
 .score_2 (score_2_x671),
 .score_3 (score_3_x671),
 .score_4 (score_4_x671),
 .score_5 (score_5_x671),
 .score_6 (score_6_x671),
 .score_7 (score_7_x671),
 .score_8 (score_8_x671),
 .score_9 (score_9_x671)
);
 
myram_28X28 #(
.ID(672),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x672),
.W_1(W_1_x672),
.W_2(W_2_x672),
.W_3(W_3_x672),
.W_4(W_4_x672),
.W_5(W_5_x672),
.W_6(W_6_x672),
.W_7(W_7_x672),
.W_8(W_8_x672),
.W_9(W_9_x672)
) u_28X28_x672 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x672),
 .score_0 (score_0_x672),
 .score_1 (score_1_x672),
 .score_2 (score_2_x672),
 .score_3 (score_3_x672),
 .score_4 (score_4_x672),
 .score_5 (score_5_x672),
 .score_6 (score_6_x672),
 .score_7 (score_7_x672),
 .score_8 (score_8_x672),
 .score_9 (score_9_x672)
);
 
myram_28X28 #(
.ID(673),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x673),
.W_1(W_1_x673),
.W_2(W_2_x673),
.W_3(W_3_x673),
.W_4(W_4_x673),
.W_5(W_5_x673),
.W_6(W_6_x673),
.W_7(W_7_x673),
.W_8(W_8_x673),
.W_9(W_9_x673)
) u_28X28_x673 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x673),
 .score_0 (score_0_x673),
 .score_1 (score_1_x673),
 .score_2 (score_2_x673),
 .score_3 (score_3_x673),
 .score_4 (score_4_x673),
 .score_5 (score_5_x673),
 .score_6 (score_6_x673),
 .score_7 (score_7_x673),
 .score_8 (score_8_x673),
 .score_9 (score_9_x673)
);
 
myram_28X28 #(
.ID(674),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x674),
.W_1(W_1_x674),
.W_2(W_2_x674),
.W_3(W_3_x674),
.W_4(W_4_x674),
.W_5(W_5_x674),
.W_6(W_6_x674),
.W_7(W_7_x674),
.W_8(W_8_x674),
.W_9(W_9_x674)
) u_28X28_x674 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x674),
 .score_0 (score_0_x674),
 .score_1 (score_1_x674),
 .score_2 (score_2_x674),
 .score_3 (score_3_x674),
 .score_4 (score_4_x674),
 .score_5 (score_5_x674),
 .score_6 (score_6_x674),
 .score_7 (score_7_x674),
 .score_8 (score_8_x674),
 .score_9 (score_9_x674)
);
 
myram_28X28 #(
.ID(675),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x675),
.W_1(W_1_x675),
.W_2(W_2_x675),
.W_3(W_3_x675),
.W_4(W_4_x675),
.W_5(W_5_x675),
.W_6(W_6_x675),
.W_7(W_7_x675),
.W_8(W_8_x675),
.W_9(W_9_x675)
) u_28X28_x675 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x675),
 .score_0 (score_0_x675),
 .score_1 (score_1_x675),
 .score_2 (score_2_x675),
 .score_3 (score_3_x675),
 .score_4 (score_4_x675),
 .score_5 (score_5_x675),
 .score_6 (score_6_x675),
 .score_7 (score_7_x675),
 .score_8 (score_8_x675),
 .score_9 (score_9_x675)
);
 
myram_28X28 #(
.ID(676),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x676),
.W_1(W_1_x676),
.W_2(W_2_x676),
.W_3(W_3_x676),
.W_4(W_4_x676),
.W_5(W_5_x676),
.W_6(W_6_x676),
.W_7(W_7_x676),
.W_8(W_8_x676),
.W_9(W_9_x676)
) u_28X28_x676 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x676),
 .score_0 (score_0_x676),
 .score_1 (score_1_x676),
 .score_2 (score_2_x676),
 .score_3 (score_3_x676),
 .score_4 (score_4_x676),
 .score_5 (score_5_x676),
 .score_6 (score_6_x676),
 .score_7 (score_7_x676),
 .score_8 (score_8_x676),
 .score_9 (score_9_x676)
);
 
myram_28X28 #(
.ID(677),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x677),
.W_1(W_1_x677),
.W_2(W_2_x677),
.W_3(W_3_x677),
.W_4(W_4_x677),
.W_5(W_5_x677),
.W_6(W_6_x677),
.W_7(W_7_x677),
.W_8(W_8_x677),
.W_9(W_9_x677)
) u_28X28_x677 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x677),
 .score_0 (score_0_x677),
 .score_1 (score_1_x677),
 .score_2 (score_2_x677),
 .score_3 (score_3_x677),
 .score_4 (score_4_x677),
 .score_5 (score_5_x677),
 .score_6 (score_6_x677),
 .score_7 (score_7_x677),
 .score_8 (score_8_x677),
 .score_9 (score_9_x677)
);
 
myram_28X28 #(
.ID(678),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x678),
.W_1(W_1_x678),
.W_2(W_2_x678),
.W_3(W_3_x678),
.W_4(W_4_x678),
.W_5(W_5_x678),
.W_6(W_6_x678),
.W_7(W_7_x678),
.W_8(W_8_x678),
.W_9(W_9_x678)
) u_28X28_x678 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x678),
 .score_0 (score_0_x678),
 .score_1 (score_1_x678),
 .score_2 (score_2_x678),
 .score_3 (score_3_x678),
 .score_4 (score_4_x678),
 .score_5 (score_5_x678),
 .score_6 (score_6_x678),
 .score_7 (score_7_x678),
 .score_8 (score_8_x678),
 .score_9 (score_9_x678)
);
 
myram_28X28 #(
.ID(679),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x679),
.W_1(W_1_x679),
.W_2(W_2_x679),
.W_3(W_3_x679),
.W_4(W_4_x679),
.W_5(W_5_x679),
.W_6(W_6_x679),
.W_7(W_7_x679),
.W_8(W_8_x679),
.W_9(W_9_x679)
) u_28X28_x679 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x679),
 .score_0 (score_0_x679),
 .score_1 (score_1_x679),
 .score_2 (score_2_x679),
 .score_3 (score_3_x679),
 .score_4 (score_4_x679),
 .score_5 (score_5_x679),
 .score_6 (score_6_x679),
 .score_7 (score_7_x679),
 .score_8 (score_8_x679),
 .score_9 (score_9_x679)
);
 
myram_28X28 #(
.ID(680),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x680),
.W_1(W_1_x680),
.W_2(W_2_x680),
.W_3(W_3_x680),
.W_4(W_4_x680),
.W_5(W_5_x680),
.W_6(W_6_x680),
.W_7(W_7_x680),
.W_8(W_8_x680),
.W_9(W_9_x680)
) u_28X28_x680 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x680),
 .score_0 (score_0_x680),
 .score_1 (score_1_x680),
 .score_2 (score_2_x680),
 .score_3 (score_3_x680),
 .score_4 (score_4_x680),
 .score_5 (score_5_x680),
 .score_6 (score_6_x680),
 .score_7 (score_7_x680),
 .score_8 (score_8_x680),
 .score_9 (score_9_x680)
);
 
myram_28X28 #(
.ID(681),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x681),
.W_1(W_1_x681),
.W_2(W_2_x681),
.W_3(W_3_x681),
.W_4(W_4_x681),
.W_5(W_5_x681),
.W_6(W_6_x681),
.W_7(W_7_x681),
.W_8(W_8_x681),
.W_9(W_9_x681)
) u_28X28_x681 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x681),
 .score_0 (score_0_x681),
 .score_1 (score_1_x681),
 .score_2 (score_2_x681),
 .score_3 (score_3_x681),
 .score_4 (score_4_x681),
 .score_5 (score_5_x681),
 .score_6 (score_6_x681),
 .score_7 (score_7_x681),
 .score_8 (score_8_x681),
 .score_9 (score_9_x681)
);
 
myram_28X28 #(
.ID(682),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x682),
.W_1(W_1_x682),
.W_2(W_2_x682),
.W_3(W_3_x682),
.W_4(W_4_x682),
.W_5(W_5_x682),
.W_6(W_6_x682),
.W_7(W_7_x682),
.W_8(W_8_x682),
.W_9(W_9_x682)
) u_28X28_x682 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x682),
 .score_0 (score_0_x682),
 .score_1 (score_1_x682),
 .score_2 (score_2_x682),
 .score_3 (score_3_x682),
 .score_4 (score_4_x682),
 .score_5 (score_5_x682),
 .score_6 (score_6_x682),
 .score_7 (score_7_x682),
 .score_8 (score_8_x682),
 .score_9 (score_9_x682)
);
 
myram_28X28 #(
.ID(683),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x683),
.W_1(W_1_x683),
.W_2(W_2_x683),
.W_3(W_3_x683),
.W_4(W_4_x683),
.W_5(W_5_x683),
.W_6(W_6_x683),
.W_7(W_7_x683),
.W_8(W_8_x683),
.W_9(W_9_x683)
) u_28X28_x683 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x683),
 .score_0 (score_0_x683),
 .score_1 (score_1_x683),
 .score_2 (score_2_x683),
 .score_3 (score_3_x683),
 .score_4 (score_4_x683),
 .score_5 (score_5_x683),
 .score_6 (score_6_x683),
 .score_7 (score_7_x683),
 .score_8 (score_8_x683),
 .score_9 (score_9_x683)
);
 
myram_28X28 #(
.ID(684),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x684),
.W_1(W_1_x684),
.W_2(W_2_x684),
.W_3(W_3_x684),
.W_4(W_4_x684),
.W_5(W_5_x684),
.W_6(W_6_x684),
.W_7(W_7_x684),
.W_8(W_8_x684),
.W_9(W_9_x684)
) u_28X28_x684 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x684),
 .score_0 (score_0_x684),
 .score_1 (score_1_x684),
 .score_2 (score_2_x684),
 .score_3 (score_3_x684),
 .score_4 (score_4_x684),
 .score_5 (score_5_x684),
 .score_6 (score_6_x684),
 .score_7 (score_7_x684),
 .score_8 (score_8_x684),
 .score_9 (score_9_x684)
);
 
myram_28X28 #(
.ID(685),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x685),
.W_1(W_1_x685),
.W_2(W_2_x685),
.W_3(W_3_x685),
.W_4(W_4_x685),
.W_5(W_5_x685),
.W_6(W_6_x685),
.W_7(W_7_x685),
.W_8(W_8_x685),
.W_9(W_9_x685)
) u_28X28_x685 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x685),
 .score_0 (score_0_x685),
 .score_1 (score_1_x685),
 .score_2 (score_2_x685),
 .score_3 (score_3_x685),
 .score_4 (score_4_x685),
 .score_5 (score_5_x685),
 .score_6 (score_6_x685),
 .score_7 (score_7_x685),
 .score_8 (score_8_x685),
 .score_9 (score_9_x685)
);
 
myram_28X28 #(
.ID(686),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x686),
.W_1(W_1_x686),
.W_2(W_2_x686),
.W_3(W_3_x686),
.W_4(W_4_x686),
.W_5(W_5_x686),
.W_6(W_6_x686),
.W_7(W_7_x686),
.W_8(W_8_x686),
.W_9(W_9_x686)
) u_28X28_x686 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x686),
 .score_0 (score_0_x686),
 .score_1 (score_1_x686),
 .score_2 (score_2_x686),
 .score_3 (score_3_x686),
 .score_4 (score_4_x686),
 .score_5 (score_5_x686),
 .score_6 (score_6_x686),
 .score_7 (score_7_x686),
 .score_8 (score_8_x686),
 .score_9 (score_9_x686)
);
 
myram_28X28 #(
.ID(687),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x687),
.W_1(W_1_x687),
.W_2(W_2_x687),
.W_3(W_3_x687),
.W_4(W_4_x687),
.W_5(W_5_x687),
.W_6(W_6_x687),
.W_7(W_7_x687),
.W_8(W_8_x687),
.W_9(W_9_x687)
) u_28X28_x687 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x687),
 .score_0 (score_0_x687),
 .score_1 (score_1_x687),
 .score_2 (score_2_x687),
 .score_3 (score_3_x687),
 .score_4 (score_4_x687),
 .score_5 (score_5_x687),
 .score_6 (score_6_x687),
 .score_7 (score_7_x687),
 .score_8 (score_8_x687),
 .score_9 (score_9_x687)
);
 
myram_28X28 #(
.ID(688),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x688),
.W_1(W_1_x688),
.W_2(W_2_x688),
.W_3(W_3_x688),
.W_4(W_4_x688),
.W_5(W_5_x688),
.W_6(W_6_x688),
.W_7(W_7_x688),
.W_8(W_8_x688),
.W_9(W_9_x688)
) u_28X28_x688 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x688),
 .score_0 (score_0_x688),
 .score_1 (score_1_x688),
 .score_2 (score_2_x688),
 .score_3 (score_3_x688),
 .score_4 (score_4_x688),
 .score_5 (score_5_x688),
 .score_6 (score_6_x688),
 .score_7 (score_7_x688),
 .score_8 (score_8_x688),
 .score_9 (score_9_x688)
);
 
myram_28X28 #(
.ID(689),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x689),
.W_1(W_1_x689),
.W_2(W_2_x689),
.W_3(W_3_x689),
.W_4(W_4_x689),
.W_5(W_5_x689),
.W_6(W_6_x689),
.W_7(W_7_x689),
.W_8(W_8_x689),
.W_9(W_9_x689)
) u_28X28_x689 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x689),
 .score_0 (score_0_x689),
 .score_1 (score_1_x689),
 .score_2 (score_2_x689),
 .score_3 (score_3_x689),
 .score_4 (score_4_x689),
 .score_5 (score_5_x689),
 .score_6 (score_6_x689),
 .score_7 (score_7_x689),
 .score_8 (score_8_x689),
 .score_9 (score_9_x689)
);
 
myram_28X28 #(
.ID(690),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x690),
.W_1(W_1_x690),
.W_2(W_2_x690),
.W_3(W_3_x690),
.W_4(W_4_x690),
.W_5(W_5_x690),
.W_6(W_6_x690),
.W_7(W_7_x690),
.W_8(W_8_x690),
.W_9(W_9_x690)
) u_28X28_x690 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x690),
 .score_0 (score_0_x690),
 .score_1 (score_1_x690),
 .score_2 (score_2_x690),
 .score_3 (score_3_x690),
 .score_4 (score_4_x690),
 .score_5 (score_5_x690),
 .score_6 (score_6_x690),
 .score_7 (score_7_x690),
 .score_8 (score_8_x690),
 .score_9 (score_9_x690)
);
 
myram_28X28 #(
.ID(691),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x691),
.W_1(W_1_x691),
.W_2(W_2_x691),
.W_3(W_3_x691),
.W_4(W_4_x691),
.W_5(W_5_x691),
.W_6(W_6_x691),
.W_7(W_7_x691),
.W_8(W_8_x691),
.W_9(W_9_x691)
) u_28X28_x691 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x691),
 .score_0 (score_0_x691),
 .score_1 (score_1_x691),
 .score_2 (score_2_x691),
 .score_3 (score_3_x691),
 .score_4 (score_4_x691),
 .score_5 (score_5_x691),
 .score_6 (score_6_x691),
 .score_7 (score_7_x691),
 .score_8 (score_8_x691),
 .score_9 (score_9_x691)
);
 
myram_28X28 #(
.ID(692),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x692),
.W_1(W_1_x692),
.W_2(W_2_x692),
.W_3(W_3_x692),
.W_4(W_4_x692),
.W_5(W_5_x692),
.W_6(W_6_x692),
.W_7(W_7_x692),
.W_8(W_8_x692),
.W_9(W_9_x692)
) u_28X28_x692 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x692),
 .score_0 (score_0_x692),
 .score_1 (score_1_x692),
 .score_2 (score_2_x692),
 .score_3 (score_3_x692),
 .score_4 (score_4_x692),
 .score_5 (score_5_x692),
 .score_6 (score_6_x692),
 .score_7 (score_7_x692),
 .score_8 (score_8_x692),
 .score_9 (score_9_x692)
);
 
myram_28X28 #(
.ID(693),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x693),
.W_1(W_1_x693),
.W_2(W_2_x693),
.W_3(W_3_x693),
.W_4(W_4_x693),
.W_5(W_5_x693),
.W_6(W_6_x693),
.W_7(W_7_x693),
.W_8(W_8_x693),
.W_9(W_9_x693)
) u_28X28_x693 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x693),
 .score_0 (score_0_x693),
 .score_1 (score_1_x693),
 .score_2 (score_2_x693),
 .score_3 (score_3_x693),
 .score_4 (score_4_x693),
 .score_5 (score_5_x693),
 .score_6 (score_6_x693),
 .score_7 (score_7_x693),
 .score_8 (score_8_x693),
 .score_9 (score_9_x693)
);
 
myram_28X28 #(
.ID(694),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x694),
.W_1(W_1_x694),
.W_2(W_2_x694),
.W_3(W_3_x694),
.W_4(W_4_x694),
.W_5(W_5_x694),
.W_6(W_6_x694),
.W_7(W_7_x694),
.W_8(W_8_x694),
.W_9(W_9_x694)
) u_28X28_x694 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x694),
 .score_0 (score_0_x694),
 .score_1 (score_1_x694),
 .score_2 (score_2_x694),
 .score_3 (score_3_x694),
 .score_4 (score_4_x694),
 .score_5 (score_5_x694),
 .score_6 (score_6_x694),
 .score_7 (score_7_x694),
 .score_8 (score_8_x694),
 .score_9 (score_9_x694)
);
 
myram_28X28 #(
.ID(695),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x695),
.W_1(W_1_x695),
.W_2(W_2_x695),
.W_3(W_3_x695),
.W_4(W_4_x695),
.W_5(W_5_x695),
.W_6(W_6_x695),
.W_7(W_7_x695),
.W_8(W_8_x695),
.W_9(W_9_x695)
) u_28X28_x695 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x695),
 .score_0 (score_0_x695),
 .score_1 (score_1_x695),
 .score_2 (score_2_x695),
 .score_3 (score_3_x695),
 .score_4 (score_4_x695),
 .score_5 (score_5_x695),
 .score_6 (score_6_x695),
 .score_7 (score_7_x695),
 .score_8 (score_8_x695),
 .score_9 (score_9_x695)
);
 
myram_28X28 #(
.ID(696),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x696),
.W_1(W_1_x696),
.W_2(W_2_x696),
.W_3(W_3_x696),
.W_4(W_4_x696),
.W_5(W_5_x696),
.W_6(W_6_x696),
.W_7(W_7_x696),
.W_8(W_8_x696),
.W_9(W_9_x696)
) u_28X28_x696 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x696),
 .score_0 (score_0_x696),
 .score_1 (score_1_x696),
 .score_2 (score_2_x696),
 .score_3 (score_3_x696),
 .score_4 (score_4_x696),
 .score_5 (score_5_x696),
 .score_6 (score_6_x696),
 .score_7 (score_7_x696),
 .score_8 (score_8_x696),
 .score_9 (score_9_x696)
);
 
myram_28X28 #(
.ID(697),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x697),
.W_1(W_1_x697),
.W_2(W_2_x697),
.W_3(W_3_x697),
.W_4(W_4_x697),
.W_5(W_5_x697),
.W_6(W_6_x697),
.W_7(W_7_x697),
.W_8(W_8_x697),
.W_9(W_9_x697)
) u_28X28_x697 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x697),
 .score_0 (score_0_x697),
 .score_1 (score_1_x697),
 .score_2 (score_2_x697),
 .score_3 (score_3_x697),
 .score_4 (score_4_x697),
 .score_5 (score_5_x697),
 .score_6 (score_6_x697),
 .score_7 (score_7_x697),
 .score_8 (score_8_x697),
 .score_9 (score_9_x697)
);
 
myram_28X28 #(
.ID(698),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x698),
.W_1(W_1_x698),
.W_2(W_2_x698),
.W_3(W_3_x698),
.W_4(W_4_x698),
.W_5(W_5_x698),
.W_6(W_6_x698),
.W_7(W_7_x698),
.W_8(W_8_x698),
.W_9(W_9_x698)
) u_28X28_x698 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x698),
 .score_0 (score_0_x698),
 .score_1 (score_1_x698),
 .score_2 (score_2_x698),
 .score_3 (score_3_x698),
 .score_4 (score_4_x698),
 .score_5 (score_5_x698),
 .score_6 (score_6_x698),
 .score_7 (score_7_x698),
 .score_8 (score_8_x698),
 .score_9 (score_9_x698)
);
 
myram_28X28 #(
.ID(699),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x699),
.W_1(W_1_x699),
.W_2(W_2_x699),
.W_3(W_3_x699),
.W_4(W_4_x699),
.W_5(W_5_x699),
.W_6(W_6_x699),
.W_7(W_7_x699),
.W_8(W_8_x699),
.W_9(W_9_x699)
) u_28X28_x699 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x699),
 .score_0 (score_0_x699),
 .score_1 (score_1_x699),
 .score_2 (score_2_x699),
 .score_3 (score_3_x699),
 .score_4 (score_4_x699),
 .score_5 (score_5_x699),
 .score_6 (score_6_x699),
 .score_7 (score_7_x699),
 .score_8 (score_8_x699),
 .score_9 (score_9_x699)
);
 
myram_28X28 #(
.ID(700),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x700),
.W_1(W_1_x700),
.W_2(W_2_x700),
.W_3(W_3_x700),
.W_4(W_4_x700),
.W_5(W_5_x700),
.W_6(W_6_x700),
.W_7(W_7_x700),
.W_8(W_8_x700),
.W_9(W_9_x700)
) u_28X28_x700 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x700),
 .score_0 (score_0_x700),
 .score_1 (score_1_x700),
 .score_2 (score_2_x700),
 .score_3 (score_3_x700),
 .score_4 (score_4_x700),
 .score_5 (score_5_x700),
 .score_6 (score_6_x700),
 .score_7 (score_7_x700),
 .score_8 (score_8_x700),
 .score_9 (score_9_x700)
);
 
myram_28X28 #(
.ID(701),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x701),
.W_1(W_1_x701),
.W_2(W_2_x701),
.W_3(W_3_x701),
.W_4(W_4_x701),
.W_5(W_5_x701),
.W_6(W_6_x701),
.W_7(W_7_x701),
.W_8(W_8_x701),
.W_9(W_9_x701)
) u_28X28_x701 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x701),
 .score_0 (score_0_x701),
 .score_1 (score_1_x701),
 .score_2 (score_2_x701),
 .score_3 (score_3_x701),
 .score_4 (score_4_x701),
 .score_5 (score_5_x701),
 .score_6 (score_6_x701),
 .score_7 (score_7_x701),
 .score_8 (score_8_x701),
 .score_9 (score_9_x701)
);
 
myram_28X28 #(
.ID(702),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x702),
.W_1(W_1_x702),
.W_2(W_2_x702),
.W_3(W_3_x702),
.W_4(W_4_x702),
.W_5(W_5_x702),
.W_6(W_6_x702),
.W_7(W_7_x702),
.W_8(W_8_x702),
.W_9(W_9_x702)
) u_28X28_x702 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x702),
 .score_0 (score_0_x702),
 .score_1 (score_1_x702),
 .score_2 (score_2_x702),
 .score_3 (score_3_x702),
 .score_4 (score_4_x702),
 .score_5 (score_5_x702),
 .score_6 (score_6_x702),
 .score_7 (score_7_x702),
 .score_8 (score_8_x702),
 .score_9 (score_9_x702)
);
 
myram_28X28 #(
.ID(703),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x703),
.W_1(W_1_x703),
.W_2(W_2_x703),
.W_3(W_3_x703),
.W_4(W_4_x703),
.W_5(W_5_x703),
.W_6(W_6_x703),
.W_7(W_7_x703),
.W_8(W_8_x703),
.W_9(W_9_x703)
) u_28X28_x703 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x703),
 .score_0 (score_0_x703),
 .score_1 (score_1_x703),
 .score_2 (score_2_x703),
 .score_3 (score_3_x703),
 .score_4 (score_4_x703),
 .score_5 (score_5_x703),
 .score_6 (score_6_x703),
 .score_7 (score_7_x703),
 .score_8 (score_8_x703),
 .score_9 (score_9_x703)
);
 
myram_28X28 #(
.ID(704),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x704),
.W_1(W_1_x704),
.W_2(W_2_x704),
.W_3(W_3_x704),
.W_4(W_4_x704),
.W_5(W_5_x704),
.W_6(W_6_x704),
.W_7(W_7_x704),
.W_8(W_8_x704),
.W_9(W_9_x704)
) u_28X28_x704 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x704),
 .score_0 (score_0_x704),
 .score_1 (score_1_x704),
 .score_2 (score_2_x704),
 .score_3 (score_3_x704),
 .score_4 (score_4_x704),
 .score_5 (score_5_x704),
 .score_6 (score_6_x704),
 .score_7 (score_7_x704),
 .score_8 (score_8_x704),
 .score_9 (score_9_x704)
);
 
myram_28X28 #(
.ID(705),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x705),
.W_1(W_1_x705),
.W_2(W_2_x705),
.W_3(W_3_x705),
.W_4(W_4_x705),
.W_5(W_5_x705),
.W_6(W_6_x705),
.W_7(W_7_x705),
.W_8(W_8_x705),
.W_9(W_9_x705)
) u_28X28_x705 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x705),
 .score_0 (score_0_x705),
 .score_1 (score_1_x705),
 .score_2 (score_2_x705),
 .score_3 (score_3_x705),
 .score_4 (score_4_x705),
 .score_5 (score_5_x705),
 .score_6 (score_6_x705),
 .score_7 (score_7_x705),
 .score_8 (score_8_x705),
 .score_9 (score_9_x705)
);
 
myram_28X28 #(
.ID(706),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x706),
.W_1(W_1_x706),
.W_2(W_2_x706),
.W_3(W_3_x706),
.W_4(W_4_x706),
.W_5(W_5_x706),
.W_6(W_6_x706),
.W_7(W_7_x706),
.W_8(W_8_x706),
.W_9(W_9_x706)
) u_28X28_x706 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x706),
 .score_0 (score_0_x706),
 .score_1 (score_1_x706),
 .score_2 (score_2_x706),
 .score_3 (score_3_x706),
 .score_4 (score_4_x706),
 .score_5 (score_5_x706),
 .score_6 (score_6_x706),
 .score_7 (score_7_x706),
 .score_8 (score_8_x706),
 .score_9 (score_9_x706)
);
 
myram_28X28 #(
.ID(707),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x707),
.W_1(W_1_x707),
.W_2(W_2_x707),
.W_3(W_3_x707),
.W_4(W_4_x707),
.W_5(W_5_x707),
.W_6(W_6_x707),
.W_7(W_7_x707),
.W_8(W_8_x707),
.W_9(W_9_x707)
) u_28X28_x707 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x707),
 .score_0 (score_0_x707),
 .score_1 (score_1_x707),
 .score_2 (score_2_x707),
 .score_3 (score_3_x707),
 .score_4 (score_4_x707),
 .score_5 (score_5_x707),
 .score_6 (score_6_x707),
 .score_7 (score_7_x707),
 .score_8 (score_8_x707),
 .score_9 (score_9_x707)
);
 
myram_28X28 #(
.ID(708),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x708),
.W_1(W_1_x708),
.W_2(W_2_x708),
.W_3(W_3_x708),
.W_4(W_4_x708),
.W_5(W_5_x708),
.W_6(W_6_x708),
.W_7(W_7_x708),
.W_8(W_8_x708),
.W_9(W_9_x708)
) u_28X28_x708 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x708),
 .score_0 (score_0_x708),
 .score_1 (score_1_x708),
 .score_2 (score_2_x708),
 .score_3 (score_3_x708),
 .score_4 (score_4_x708),
 .score_5 (score_5_x708),
 .score_6 (score_6_x708),
 .score_7 (score_7_x708),
 .score_8 (score_8_x708),
 .score_9 (score_9_x708)
);
 
myram_28X28 #(
.ID(709),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x709),
.W_1(W_1_x709),
.W_2(W_2_x709),
.W_3(W_3_x709),
.W_4(W_4_x709),
.W_5(W_5_x709),
.W_6(W_6_x709),
.W_7(W_7_x709),
.W_8(W_8_x709),
.W_9(W_9_x709)
) u_28X28_x709 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x709),
 .score_0 (score_0_x709),
 .score_1 (score_1_x709),
 .score_2 (score_2_x709),
 .score_3 (score_3_x709),
 .score_4 (score_4_x709),
 .score_5 (score_5_x709),
 .score_6 (score_6_x709),
 .score_7 (score_7_x709),
 .score_8 (score_8_x709),
 .score_9 (score_9_x709)
);
 
myram_28X28 #(
.ID(710),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x710),
.W_1(W_1_x710),
.W_2(W_2_x710),
.W_3(W_3_x710),
.W_4(W_4_x710),
.W_5(W_5_x710),
.W_6(W_6_x710),
.W_7(W_7_x710),
.W_8(W_8_x710),
.W_9(W_9_x710)
) u_28X28_x710 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x710),
 .score_0 (score_0_x710),
 .score_1 (score_1_x710),
 .score_2 (score_2_x710),
 .score_3 (score_3_x710),
 .score_4 (score_4_x710),
 .score_5 (score_5_x710),
 .score_6 (score_6_x710),
 .score_7 (score_7_x710),
 .score_8 (score_8_x710),
 .score_9 (score_9_x710)
);
 
myram_28X28 #(
.ID(711),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x711),
.W_1(W_1_x711),
.W_2(W_2_x711),
.W_3(W_3_x711),
.W_4(W_4_x711),
.W_5(W_5_x711),
.W_6(W_6_x711),
.W_7(W_7_x711),
.W_8(W_8_x711),
.W_9(W_9_x711)
) u_28X28_x711 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x711),
 .score_0 (score_0_x711),
 .score_1 (score_1_x711),
 .score_2 (score_2_x711),
 .score_3 (score_3_x711),
 .score_4 (score_4_x711),
 .score_5 (score_5_x711),
 .score_6 (score_6_x711),
 .score_7 (score_7_x711),
 .score_8 (score_8_x711),
 .score_9 (score_9_x711)
);
 
myram_28X28 #(
.ID(712),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x712),
.W_1(W_1_x712),
.W_2(W_2_x712),
.W_3(W_3_x712),
.W_4(W_4_x712),
.W_5(W_5_x712),
.W_6(W_6_x712),
.W_7(W_7_x712),
.W_8(W_8_x712),
.W_9(W_9_x712)
) u_28X28_x712 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x712),
 .score_0 (score_0_x712),
 .score_1 (score_1_x712),
 .score_2 (score_2_x712),
 .score_3 (score_3_x712),
 .score_4 (score_4_x712),
 .score_5 (score_5_x712),
 .score_6 (score_6_x712),
 .score_7 (score_7_x712),
 .score_8 (score_8_x712),
 .score_9 (score_9_x712)
);
 
myram_28X28 #(
.ID(713),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x713),
.W_1(W_1_x713),
.W_2(W_2_x713),
.W_3(W_3_x713),
.W_4(W_4_x713),
.W_5(W_5_x713),
.W_6(W_6_x713),
.W_7(W_7_x713),
.W_8(W_8_x713),
.W_9(W_9_x713)
) u_28X28_x713 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x713),
 .score_0 (score_0_x713),
 .score_1 (score_1_x713),
 .score_2 (score_2_x713),
 .score_3 (score_3_x713),
 .score_4 (score_4_x713),
 .score_5 (score_5_x713),
 .score_6 (score_6_x713),
 .score_7 (score_7_x713),
 .score_8 (score_8_x713),
 .score_9 (score_9_x713)
);
 
myram_28X28 #(
.ID(714),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x714),
.W_1(W_1_x714),
.W_2(W_2_x714),
.W_3(W_3_x714),
.W_4(W_4_x714),
.W_5(W_5_x714),
.W_6(W_6_x714),
.W_7(W_7_x714),
.W_8(W_8_x714),
.W_9(W_9_x714)
) u_28X28_x714 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x714),
 .score_0 (score_0_x714),
 .score_1 (score_1_x714),
 .score_2 (score_2_x714),
 .score_3 (score_3_x714),
 .score_4 (score_4_x714),
 .score_5 (score_5_x714),
 .score_6 (score_6_x714),
 .score_7 (score_7_x714),
 .score_8 (score_8_x714),
 .score_9 (score_9_x714)
);
 
myram_28X28 #(
.ID(715),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x715),
.W_1(W_1_x715),
.W_2(W_2_x715),
.W_3(W_3_x715),
.W_4(W_4_x715),
.W_5(W_5_x715),
.W_6(W_6_x715),
.W_7(W_7_x715),
.W_8(W_8_x715),
.W_9(W_9_x715)
) u_28X28_x715 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x715),
 .score_0 (score_0_x715),
 .score_1 (score_1_x715),
 .score_2 (score_2_x715),
 .score_3 (score_3_x715),
 .score_4 (score_4_x715),
 .score_5 (score_5_x715),
 .score_6 (score_6_x715),
 .score_7 (score_7_x715),
 .score_8 (score_8_x715),
 .score_9 (score_9_x715)
);
 
myram_28X28 #(
.ID(716),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x716),
.W_1(W_1_x716),
.W_2(W_2_x716),
.W_3(W_3_x716),
.W_4(W_4_x716),
.W_5(W_5_x716),
.W_6(W_6_x716),
.W_7(W_7_x716),
.W_8(W_8_x716),
.W_9(W_9_x716)
) u_28X28_x716 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x716),
 .score_0 (score_0_x716),
 .score_1 (score_1_x716),
 .score_2 (score_2_x716),
 .score_3 (score_3_x716),
 .score_4 (score_4_x716),
 .score_5 (score_5_x716),
 .score_6 (score_6_x716),
 .score_7 (score_7_x716),
 .score_8 (score_8_x716),
 .score_9 (score_9_x716)
);
 
myram_28X28 #(
.ID(717),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x717),
.W_1(W_1_x717),
.W_2(W_2_x717),
.W_3(W_3_x717),
.W_4(W_4_x717),
.W_5(W_5_x717),
.W_6(W_6_x717),
.W_7(W_7_x717),
.W_8(W_8_x717),
.W_9(W_9_x717)
) u_28X28_x717 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x717),
 .score_0 (score_0_x717),
 .score_1 (score_1_x717),
 .score_2 (score_2_x717),
 .score_3 (score_3_x717),
 .score_4 (score_4_x717),
 .score_5 (score_5_x717),
 .score_6 (score_6_x717),
 .score_7 (score_7_x717),
 .score_8 (score_8_x717),
 .score_9 (score_9_x717)
);
 
myram_28X28 #(
.ID(718),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x718),
.W_1(W_1_x718),
.W_2(W_2_x718),
.W_3(W_3_x718),
.W_4(W_4_x718),
.W_5(W_5_x718),
.W_6(W_6_x718),
.W_7(W_7_x718),
.W_8(W_8_x718),
.W_9(W_9_x718)
) u_28X28_x718 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x718),
 .score_0 (score_0_x718),
 .score_1 (score_1_x718),
 .score_2 (score_2_x718),
 .score_3 (score_3_x718),
 .score_4 (score_4_x718),
 .score_5 (score_5_x718),
 .score_6 (score_6_x718),
 .score_7 (score_7_x718),
 .score_8 (score_8_x718),
 .score_9 (score_9_x718)
);
 
myram_28X28 #(
.ID(719),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x719),
.W_1(W_1_x719),
.W_2(W_2_x719),
.W_3(W_3_x719),
.W_4(W_4_x719),
.W_5(W_5_x719),
.W_6(W_6_x719),
.W_7(W_7_x719),
.W_8(W_8_x719),
.W_9(W_9_x719)
) u_28X28_x719 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x719),
 .score_0 (score_0_x719),
 .score_1 (score_1_x719),
 .score_2 (score_2_x719),
 .score_3 (score_3_x719),
 .score_4 (score_4_x719),
 .score_5 (score_5_x719),
 .score_6 (score_6_x719),
 .score_7 (score_7_x719),
 .score_8 (score_8_x719),
 .score_9 (score_9_x719)
);
 
myram_28X28 #(
.ID(720),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x720),
.W_1(W_1_x720),
.W_2(W_2_x720),
.W_3(W_3_x720),
.W_4(W_4_x720),
.W_5(W_5_x720),
.W_6(W_6_x720),
.W_7(W_7_x720),
.W_8(W_8_x720),
.W_9(W_9_x720)
) u_28X28_x720 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x720),
 .score_0 (score_0_x720),
 .score_1 (score_1_x720),
 .score_2 (score_2_x720),
 .score_3 (score_3_x720),
 .score_4 (score_4_x720),
 .score_5 (score_5_x720),
 .score_6 (score_6_x720),
 .score_7 (score_7_x720),
 .score_8 (score_8_x720),
 .score_9 (score_9_x720)
);
 
myram_28X28 #(
.ID(721),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x721),
.W_1(W_1_x721),
.W_2(W_2_x721),
.W_3(W_3_x721),
.W_4(W_4_x721),
.W_5(W_5_x721),
.W_6(W_6_x721),
.W_7(W_7_x721),
.W_8(W_8_x721),
.W_9(W_9_x721)
) u_28X28_x721 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x721),
 .score_0 (score_0_x721),
 .score_1 (score_1_x721),
 .score_2 (score_2_x721),
 .score_3 (score_3_x721),
 .score_4 (score_4_x721),
 .score_5 (score_5_x721),
 .score_6 (score_6_x721),
 .score_7 (score_7_x721),
 .score_8 (score_8_x721),
 .score_9 (score_9_x721)
);
 
myram_28X28 #(
.ID(722),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x722),
.W_1(W_1_x722),
.W_2(W_2_x722),
.W_3(W_3_x722),
.W_4(W_4_x722),
.W_5(W_5_x722),
.W_6(W_6_x722),
.W_7(W_7_x722),
.W_8(W_8_x722),
.W_9(W_9_x722)
) u_28X28_x722 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x722),
 .score_0 (score_0_x722),
 .score_1 (score_1_x722),
 .score_2 (score_2_x722),
 .score_3 (score_3_x722),
 .score_4 (score_4_x722),
 .score_5 (score_5_x722),
 .score_6 (score_6_x722),
 .score_7 (score_7_x722),
 .score_8 (score_8_x722),
 .score_9 (score_9_x722)
);
 
myram_28X28 #(
.ID(723),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x723),
.W_1(W_1_x723),
.W_2(W_2_x723),
.W_3(W_3_x723),
.W_4(W_4_x723),
.W_5(W_5_x723),
.W_6(W_6_x723),
.W_7(W_7_x723),
.W_8(W_8_x723),
.W_9(W_9_x723)
) u_28X28_x723 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x723),
 .score_0 (score_0_x723),
 .score_1 (score_1_x723),
 .score_2 (score_2_x723),
 .score_3 (score_3_x723),
 .score_4 (score_4_x723),
 .score_5 (score_5_x723),
 .score_6 (score_6_x723),
 .score_7 (score_7_x723),
 .score_8 (score_8_x723),
 .score_9 (score_9_x723)
);
 
myram_28X28 #(
.ID(724),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x724),
.W_1(W_1_x724),
.W_2(W_2_x724),
.W_3(W_3_x724),
.W_4(W_4_x724),
.W_5(W_5_x724),
.W_6(W_6_x724),
.W_7(W_7_x724),
.W_8(W_8_x724),
.W_9(W_9_x724)
) u_28X28_x724 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x724),
 .score_0 (score_0_x724),
 .score_1 (score_1_x724),
 .score_2 (score_2_x724),
 .score_3 (score_3_x724),
 .score_4 (score_4_x724),
 .score_5 (score_5_x724),
 .score_6 (score_6_x724),
 .score_7 (score_7_x724),
 .score_8 (score_8_x724),
 .score_9 (score_9_x724)
);
 
myram_28X28 #(
.ID(725),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x725),
.W_1(W_1_x725),
.W_2(W_2_x725),
.W_3(W_3_x725),
.W_4(W_4_x725),
.W_5(W_5_x725),
.W_6(W_6_x725),
.W_7(W_7_x725),
.W_8(W_8_x725),
.W_9(W_9_x725)
) u_28X28_x725 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x725),
 .score_0 (score_0_x725),
 .score_1 (score_1_x725),
 .score_2 (score_2_x725),
 .score_3 (score_3_x725),
 .score_4 (score_4_x725),
 .score_5 (score_5_x725),
 .score_6 (score_6_x725),
 .score_7 (score_7_x725),
 .score_8 (score_8_x725),
 .score_9 (score_9_x725)
);
 
myram_28X28 #(
.ID(726),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x726),
.W_1(W_1_x726),
.W_2(W_2_x726),
.W_3(W_3_x726),
.W_4(W_4_x726),
.W_5(W_5_x726),
.W_6(W_6_x726),
.W_7(W_7_x726),
.W_8(W_8_x726),
.W_9(W_9_x726)
) u_28X28_x726 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x726),
 .score_0 (score_0_x726),
 .score_1 (score_1_x726),
 .score_2 (score_2_x726),
 .score_3 (score_3_x726),
 .score_4 (score_4_x726),
 .score_5 (score_5_x726),
 .score_6 (score_6_x726),
 .score_7 (score_7_x726),
 .score_8 (score_8_x726),
 .score_9 (score_9_x726)
);
 
myram_28X28 #(
.ID(727),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x727),
.W_1(W_1_x727),
.W_2(W_2_x727),
.W_3(W_3_x727),
.W_4(W_4_x727),
.W_5(W_5_x727),
.W_6(W_6_x727),
.W_7(W_7_x727),
.W_8(W_8_x727),
.W_9(W_9_x727)
) u_28X28_x727 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x727),
 .score_0 (score_0_x727),
 .score_1 (score_1_x727),
 .score_2 (score_2_x727),
 .score_3 (score_3_x727),
 .score_4 (score_4_x727),
 .score_5 (score_5_x727),
 .score_6 (score_6_x727),
 .score_7 (score_7_x727),
 .score_8 (score_8_x727),
 .score_9 (score_9_x727)
);
 
myram_28X28 #(
.ID(728),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x728),
.W_1(W_1_x728),
.W_2(W_2_x728),
.W_3(W_3_x728),
.W_4(W_4_x728),
.W_5(W_5_x728),
.W_6(W_6_x728),
.W_7(W_7_x728),
.W_8(W_8_x728),
.W_9(W_9_x728)
) u_28X28_x728 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x728),
 .score_0 (score_0_x728),
 .score_1 (score_1_x728),
 .score_2 (score_2_x728),
 .score_3 (score_3_x728),
 .score_4 (score_4_x728),
 .score_5 (score_5_x728),
 .score_6 (score_6_x728),
 .score_7 (score_7_x728),
 .score_8 (score_8_x728),
 .score_9 (score_9_x728)
);
 
myram_28X28 #(
.ID(729),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x729),
.W_1(W_1_x729),
.W_2(W_2_x729),
.W_3(W_3_x729),
.W_4(W_4_x729),
.W_5(W_5_x729),
.W_6(W_6_x729),
.W_7(W_7_x729),
.W_8(W_8_x729),
.W_9(W_9_x729)
) u_28X28_x729 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x729),
 .score_0 (score_0_x729),
 .score_1 (score_1_x729),
 .score_2 (score_2_x729),
 .score_3 (score_3_x729),
 .score_4 (score_4_x729),
 .score_5 (score_5_x729),
 .score_6 (score_6_x729),
 .score_7 (score_7_x729),
 .score_8 (score_8_x729),
 .score_9 (score_9_x729)
);
 
myram_28X28 #(
.ID(730),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x730),
.W_1(W_1_x730),
.W_2(W_2_x730),
.W_3(W_3_x730),
.W_4(W_4_x730),
.W_5(W_5_x730),
.W_6(W_6_x730),
.W_7(W_7_x730),
.W_8(W_8_x730),
.W_9(W_9_x730)
) u_28X28_x730 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x730),
 .score_0 (score_0_x730),
 .score_1 (score_1_x730),
 .score_2 (score_2_x730),
 .score_3 (score_3_x730),
 .score_4 (score_4_x730),
 .score_5 (score_5_x730),
 .score_6 (score_6_x730),
 .score_7 (score_7_x730),
 .score_8 (score_8_x730),
 .score_9 (score_9_x730)
);
 
myram_28X28 #(
.ID(731),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x731),
.W_1(W_1_x731),
.W_2(W_2_x731),
.W_3(W_3_x731),
.W_4(W_4_x731),
.W_5(W_5_x731),
.W_6(W_6_x731),
.W_7(W_7_x731),
.W_8(W_8_x731),
.W_9(W_9_x731)
) u_28X28_x731 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x731),
 .score_0 (score_0_x731),
 .score_1 (score_1_x731),
 .score_2 (score_2_x731),
 .score_3 (score_3_x731),
 .score_4 (score_4_x731),
 .score_5 (score_5_x731),
 .score_6 (score_6_x731),
 .score_7 (score_7_x731),
 .score_8 (score_8_x731),
 .score_9 (score_9_x731)
);
 
myram_28X28 #(
.ID(732),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x732),
.W_1(W_1_x732),
.W_2(W_2_x732),
.W_3(W_3_x732),
.W_4(W_4_x732),
.W_5(W_5_x732),
.W_6(W_6_x732),
.W_7(W_7_x732),
.W_8(W_8_x732),
.W_9(W_9_x732)
) u_28X28_x732 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x732),
 .score_0 (score_0_x732),
 .score_1 (score_1_x732),
 .score_2 (score_2_x732),
 .score_3 (score_3_x732),
 .score_4 (score_4_x732),
 .score_5 (score_5_x732),
 .score_6 (score_6_x732),
 .score_7 (score_7_x732),
 .score_8 (score_8_x732),
 .score_9 (score_9_x732)
);
 
myram_28X28 #(
.ID(733),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x733),
.W_1(W_1_x733),
.W_2(W_2_x733),
.W_3(W_3_x733),
.W_4(W_4_x733),
.W_5(W_5_x733),
.W_6(W_6_x733),
.W_7(W_7_x733),
.W_8(W_8_x733),
.W_9(W_9_x733)
) u_28X28_x733 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x733),
 .score_0 (score_0_x733),
 .score_1 (score_1_x733),
 .score_2 (score_2_x733),
 .score_3 (score_3_x733),
 .score_4 (score_4_x733),
 .score_5 (score_5_x733),
 .score_6 (score_6_x733),
 .score_7 (score_7_x733),
 .score_8 (score_8_x733),
 .score_9 (score_9_x733)
);
 
myram_28X28 #(
.ID(734),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x734),
.W_1(W_1_x734),
.W_2(W_2_x734),
.W_3(W_3_x734),
.W_4(W_4_x734),
.W_5(W_5_x734),
.W_6(W_6_x734),
.W_7(W_7_x734),
.W_8(W_8_x734),
.W_9(W_9_x734)
) u_28X28_x734 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x734),
 .score_0 (score_0_x734),
 .score_1 (score_1_x734),
 .score_2 (score_2_x734),
 .score_3 (score_3_x734),
 .score_4 (score_4_x734),
 .score_5 (score_5_x734),
 .score_6 (score_6_x734),
 .score_7 (score_7_x734),
 .score_8 (score_8_x734),
 .score_9 (score_9_x734)
);
 
myram_28X28 #(
.ID(735),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x735),
.W_1(W_1_x735),
.W_2(W_2_x735),
.W_3(W_3_x735),
.W_4(W_4_x735),
.W_5(W_5_x735),
.W_6(W_6_x735),
.W_7(W_7_x735),
.W_8(W_8_x735),
.W_9(W_9_x735)
) u_28X28_x735 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x735),
 .score_0 (score_0_x735),
 .score_1 (score_1_x735),
 .score_2 (score_2_x735),
 .score_3 (score_3_x735),
 .score_4 (score_4_x735),
 .score_5 (score_5_x735),
 .score_6 (score_6_x735),
 .score_7 (score_7_x735),
 .score_8 (score_8_x735),
 .score_9 (score_9_x735)
);
 
myram_28X28 #(
.ID(736),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x736),
.W_1(W_1_x736),
.W_2(W_2_x736),
.W_3(W_3_x736),
.W_4(W_4_x736),
.W_5(W_5_x736),
.W_6(W_6_x736),
.W_7(W_7_x736),
.W_8(W_8_x736),
.W_9(W_9_x736)
) u_28X28_x736 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x736),
 .score_0 (score_0_x736),
 .score_1 (score_1_x736),
 .score_2 (score_2_x736),
 .score_3 (score_3_x736),
 .score_4 (score_4_x736),
 .score_5 (score_5_x736),
 .score_6 (score_6_x736),
 .score_7 (score_7_x736),
 .score_8 (score_8_x736),
 .score_9 (score_9_x736)
);
 
myram_28X28 #(
.ID(737),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x737),
.W_1(W_1_x737),
.W_2(W_2_x737),
.W_3(W_3_x737),
.W_4(W_4_x737),
.W_5(W_5_x737),
.W_6(W_6_x737),
.W_7(W_7_x737),
.W_8(W_8_x737),
.W_9(W_9_x737)
) u_28X28_x737 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x737),
 .score_0 (score_0_x737),
 .score_1 (score_1_x737),
 .score_2 (score_2_x737),
 .score_3 (score_3_x737),
 .score_4 (score_4_x737),
 .score_5 (score_5_x737),
 .score_6 (score_6_x737),
 .score_7 (score_7_x737),
 .score_8 (score_8_x737),
 .score_9 (score_9_x737)
);
 
myram_28X28 #(
.ID(738),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x738),
.W_1(W_1_x738),
.W_2(W_2_x738),
.W_3(W_3_x738),
.W_4(W_4_x738),
.W_5(W_5_x738),
.W_6(W_6_x738),
.W_7(W_7_x738),
.W_8(W_8_x738),
.W_9(W_9_x738)
) u_28X28_x738 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x738),
 .score_0 (score_0_x738),
 .score_1 (score_1_x738),
 .score_2 (score_2_x738),
 .score_3 (score_3_x738),
 .score_4 (score_4_x738),
 .score_5 (score_5_x738),
 .score_6 (score_6_x738),
 .score_7 (score_7_x738),
 .score_8 (score_8_x738),
 .score_9 (score_9_x738)
);
 
myram_28X28 #(
.ID(739),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x739),
.W_1(W_1_x739),
.W_2(W_2_x739),
.W_3(W_3_x739),
.W_4(W_4_x739),
.W_5(W_5_x739),
.W_6(W_6_x739),
.W_7(W_7_x739),
.W_8(W_8_x739),
.W_9(W_9_x739)
) u_28X28_x739 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x739),
 .score_0 (score_0_x739),
 .score_1 (score_1_x739),
 .score_2 (score_2_x739),
 .score_3 (score_3_x739),
 .score_4 (score_4_x739),
 .score_5 (score_5_x739),
 .score_6 (score_6_x739),
 .score_7 (score_7_x739),
 .score_8 (score_8_x739),
 .score_9 (score_9_x739)
);
 
myram_28X28 #(
.ID(740),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x740),
.W_1(W_1_x740),
.W_2(W_2_x740),
.W_3(W_3_x740),
.W_4(W_4_x740),
.W_5(W_5_x740),
.W_6(W_6_x740),
.W_7(W_7_x740),
.W_8(W_8_x740),
.W_9(W_9_x740)
) u_28X28_x740 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x740),
 .score_0 (score_0_x740),
 .score_1 (score_1_x740),
 .score_2 (score_2_x740),
 .score_3 (score_3_x740),
 .score_4 (score_4_x740),
 .score_5 (score_5_x740),
 .score_6 (score_6_x740),
 .score_7 (score_7_x740),
 .score_8 (score_8_x740),
 .score_9 (score_9_x740)
);
 
myram_28X28 #(
.ID(741),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x741),
.W_1(W_1_x741),
.W_2(W_2_x741),
.W_3(W_3_x741),
.W_4(W_4_x741),
.W_5(W_5_x741),
.W_6(W_6_x741),
.W_7(W_7_x741),
.W_8(W_8_x741),
.W_9(W_9_x741)
) u_28X28_x741 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x741),
 .score_0 (score_0_x741),
 .score_1 (score_1_x741),
 .score_2 (score_2_x741),
 .score_3 (score_3_x741),
 .score_4 (score_4_x741),
 .score_5 (score_5_x741),
 .score_6 (score_6_x741),
 .score_7 (score_7_x741),
 .score_8 (score_8_x741),
 .score_9 (score_9_x741)
);
 
myram_28X28 #(
.ID(742),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x742),
.W_1(W_1_x742),
.W_2(W_2_x742),
.W_3(W_3_x742),
.W_4(W_4_x742),
.W_5(W_5_x742),
.W_6(W_6_x742),
.W_7(W_7_x742),
.W_8(W_8_x742),
.W_9(W_9_x742)
) u_28X28_x742 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x742),
 .score_0 (score_0_x742),
 .score_1 (score_1_x742),
 .score_2 (score_2_x742),
 .score_3 (score_3_x742),
 .score_4 (score_4_x742),
 .score_5 (score_5_x742),
 .score_6 (score_6_x742),
 .score_7 (score_7_x742),
 .score_8 (score_8_x742),
 .score_9 (score_9_x742)
);
 
myram_28X28 #(
.ID(743),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x743),
.W_1(W_1_x743),
.W_2(W_2_x743),
.W_3(W_3_x743),
.W_4(W_4_x743),
.W_5(W_5_x743),
.W_6(W_6_x743),
.W_7(W_7_x743),
.W_8(W_8_x743),
.W_9(W_9_x743)
) u_28X28_x743 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x743),
 .score_0 (score_0_x743),
 .score_1 (score_1_x743),
 .score_2 (score_2_x743),
 .score_3 (score_3_x743),
 .score_4 (score_4_x743),
 .score_5 (score_5_x743),
 .score_6 (score_6_x743),
 .score_7 (score_7_x743),
 .score_8 (score_8_x743),
 .score_9 (score_9_x743)
);
 
myram_28X28 #(
.ID(744),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x744),
.W_1(W_1_x744),
.W_2(W_2_x744),
.W_3(W_3_x744),
.W_4(W_4_x744),
.W_5(W_5_x744),
.W_6(W_6_x744),
.W_7(W_7_x744),
.W_8(W_8_x744),
.W_9(W_9_x744)
) u_28X28_x744 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x744),
 .score_0 (score_0_x744),
 .score_1 (score_1_x744),
 .score_2 (score_2_x744),
 .score_3 (score_3_x744),
 .score_4 (score_4_x744),
 .score_5 (score_5_x744),
 .score_6 (score_6_x744),
 .score_7 (score_7_x744),
 .score_8 (score_8_x744),
 .score_9 (score_9_x744)
);
 
myram_28X28 #(
.ID(745),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x745),
.W_1(W_1_x745),
.W_2(W_2_x745),
.W_3(W_3_x745),
.W_4(W_4_x745),
.W_5(W_5_x745),
.W_6(W_6_x745),
.W_7(W_7_x745),
.W_8(W_8_x745),
.W_9(W_9_x745)
) u_28X28_x745 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x745),
 .score_0 (score_0_x745),
 .score_1 (score_1_x745),
 .score_2 (score_2_x745),
 .score_3 (score_3_x745),
 .score_4 (score_4_x745),
 .score_5 (score_5_x745),
 .score_6 (score_6_x745),
 .score_7 (score_7_x745),
 .score_8 (score_8_x745),
 .score_9 (score_9_x745)
);
 
myram_28X28 #(
.ID(746),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x746),
.W_1(W_1_x746),
.W_2(W_2_x746),
.W_3(W_3_x746),
.W_4(W_4_x746),
.W_5(W_5_x746),
.W_6(W_6_x746),
.W_7(W_7_x746),
.W_8(W_8_x746),
.W_9(W_9_x746)
) u_28X28_x746 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x746),
 .score_0 (score_0_x746),
 .score_1 (score_1_x746),
 .score_2 (score_2_x746),
 .score_3 (score_3_x746),
 .score_4 (score_4_x746),
 .score_5 (score_5_x746),
 .score_6 (score_6_x746),
 .score_7 (score_7_x746),
 .score_8 (score_8_x746),
 .score_9 (score_9_x746)
);
 
myram_28X28 #(
.ID(747),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x747),
.W_1(W_1_x747),
.W_2(W_2_x747),
.W_3(W_3_x747),
.W_4(W_4_x747),
.W_5(W_5_x747),
.W_6(W_6_x747),
.W_7(W_7_x747),
.W_8(W_8_x747),
.W_9(W_9_x747)
) u_28X28_x747 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x747),
 .score_0 (score_0_x747),
 .score_1 (score_1_x747),
 .score_2 (score_2_x747),
 .score_3 (score_3_x747),
 .score_4 (score_4_x747),
 .score_5 (score_5_x747),
 .score_6 (score_6_x747),
 .score_7 (score_7_x747),
 .score_8 (score_8_x747),
 .score_9 (score_9_x747)
);
 
myram_28X28 #(
.ID(748),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x748),
.W_1(W_1_x748),
.W_2(W_2_x748),
.W_3(W_3_x748),
.W_4(W_4_x748),
.W_5(W_5_x748),
.W_6(W_6_x748),
.W_7(W_7_x748),
.W_8(W_8_x748),
.W_9(W_9_x748)
) u_28X28_x748 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x748),
 .score_0 (score_0_x748),
 .score_1 (score_1_x748),
 .score_2 (score_2_x748),
 .score_3 (score_3_x748),
 .score_4 (score_4_x748),
 .score_5 (score_5_x748),
 .score_6 (score_6_x748),
 .score_7 (score_7_x748),
 .score_8 (score_8_x748),
 .score_9 (score_9_x748)
);
 
myram_28X28 #(
.ID(749),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x749),
.W_1(W_1_x749),
.W_2(W_2_x749),
.W_3(W_3_x749),
.W_4(W_4_x749),
.W_5(W_5_x749),
.W_6(W_6_x749),
.W_7(W_7_x749),
.W_8(W_8_x749),
.W_9(W_9_x749)
) u_28X28_x749 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x749),
 .score_0 (score_0_x749),
 .score_1 (score_1_x749),
 .score_2 (score_2_x749),
 .score_3 (score_3_x749),
 .score_4 (score_4_x749),
 .score_5 (score_5_x749),
 .score_6 (score_6_x749),
 .score_7 (score_7_x749),
 .score_8 (score_8_x749),
 .score_9 (score_9_x749)
);
 
myram_28X28 #(
.ID(750),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x750),
.W_1(W_1_x750),
.W_2(W_2_x750),
.W_3(W_3_x750),
.W_4(W_4_x750),
.W_5(W_5_x750),
.W_6(W_6_x750),
.W_7(W_7_x750),
.W_8(W_8_x750),
.W_9(W_9_x750)
) u_28X28_x750 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x750),
 .score_0 (score_0_x750),
 .score_1 (score_1_x750),
 .score_2 (score_2_x750),
 .score_3 (score_3_x750),
 .score_4 (score_4_x750),
 .score_5 (score_5_x750),
 .score_6 (score_6_x750),
 .score_7 (score_7_x750),
 .score_8 (score_8_x750),
 .score_9 (score_9_x750)
);
 
myram_28X28 #(
.ID(751),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x751),
.W_1(W_1_x751),
.W_2(W_2_x751),
.W_3(W_3_x751),
.W_4(W_4_x751),
.W_5(W_5_x751),
.W_6(W_6_x751),
.W_7(W_7_x751),
.W_8(W_8_x751),
.W_9(W_9_x751)
) u_28X28_x751 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x751),
 .score_0 (score_0_x751),
 .score_1 (score_1_x751),
 .score_2 (score_2_x751),
 .score_3 (score_3_x751),
 .score_4 (score_4_x751),
 .score_5 (score_5_x751),
 .score_6 (score_6_x751),
 .score_7 (score_7_x751),
 .score_8 (score_8_x751),
 .score_9 (score_9_x751)
);
 
myram_28X28 #(
.ID(752),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x752),
.W_1(W_1_x752),
.W_2(W_2_x752),
.W_3(W_3_x752),
.W_4(W_4_x752),
.W_5(W_5_x752),
.W_6(W_6_x752),
.W_7(W_7_x752),
.W_8(W_8_x752),
.W_9(W_9_x752)
) u_28X28_x752 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x752),
 .score_0 (score_0_x752),
 .score_1 (score_1_x752),
 .score_2 (score_2_x752),
 .score_3 (score_3_x752),
 .score_4 (score_4_x752),
 .score_5 (score_5_x752),
 .score_6 (score_6_x752),
 .score_7 (score_7_x752),
 .score_8 (score_8_x752),
 .score_9 (score_9_x752)
);
 
myram_28X28 #(
.ID(753),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x753),
.W_1(W_1_x753),
.W_2(W_2_x753),
.W_3(W_3_x753),
.W_4(W_4_x753),
.W_5(W_5_x753),
.W_6(W_6_x753),
.W_7(W_7_x753),
.W_8(W_8_x753),
.W_9(W_9_x753)
) u_28X28_x753 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x753),
 .score_0 (score_0_x753),
 .score_1 (score_1_x753),
 .score_2 (score_2_x753),
 .score_3 (score_3_x753),
 .score_4 (score_4_x753),
 .score_5 (score_5_x753),
 .score_6 (score_6_x753),
 .score_7 (score_7_x753),
 .score_8 (score_8_x753),
 .score_9 (score_9_x753)
);
 
myram_28X28 #(
.ID(754),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x754),
.W_1(W_1_x754),
.W_2(W_2_x754),
.W_3(W_3_x754),
.W_4(W_4_x754),
.W_5(W_5_x754),
.W_6(W_6_x754),
.W_7(W_7_x754),
.W_8(W_8_x754),
.W_9(W_9_x754)
) u_28X28_x754 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x754),
 .score_0 (score_0_x754),
 .score_1 (score_1_x754),
 .score_2 (score_2_x754),
 .score_3 (score_3_x754),
 .score_4 (score_4_x754),
 .score_5 (score_5_x754),
 .score_6 (score_6_x754),
 .score_7 (score_7_x754),
 .score_8 (score_8_x754),
 .score_9 (score_9_x754)
);
 
myram_28X28 #(
.ID(755),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x755),
.W_1(W_1_x755),
.W_2(W_2_x755),
.W_3(W_3_x755),
.W_4(W_4_x755),
.W_5(W_5_x755),
.W_6(W_6_x755),
.W_7(W_7_x755),
.W_8(W_8_x755),
.W_9(W_9_x755)
) u_28X28_x755 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x755),
 .score_0 (score_0_x755),
 .score_1 (score_1_x755),
 .score_2 (score_2_x755),
 .score_3 (score_3_x755),
 .score_4 (score_4_x755),
 .score_5 (score_5_x755),
 .score_6 (score_6_x755),
 .score_7 (score_7_x755),
 .score_8 (score_8_x755),
 .score_9 (score_9_x755)
);
 
myram_28X28 #(
.ID(756),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x756),
.W_1(W_1_x756),
.W_2(W_2_x756),
.W_3(W_3_x756),
.W_4(W_4_x756),
.W_5(W_5_x756),
.W_6(W_6_x756),
.W_7(W_7_x756),
.W_8(W_8_x756),
.W_9(W_9_x756)
) u_28X28_x756 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x756),
 .score_0 (score_0_x756),
 .score_1 (score_1_x756),
 .score_2 (score_2_x756),
 .score_3 (score_3_x756),
 .score_4 (score_4_x756),
 .score_5 (score_5_x756),
 .score_6 (score_6_x756),
 .score_7 (score_7_x756),
 .score_8 (score_8_x756),
 .score_9 (score_9_x756)
);
 
myram_28X28 #(
.ID(757),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x757),
.W_1(W_1_x757),
.W_2(W_2_x757),
.W_3(W_3_x757),
.W_4(W_4_x757),
.W_5(W_5_x757),
.W_6(W_6_x757),
.W_7(W_7_x757),
.W_8(W_8_x757),
.W_9(W_9_x757)
) u_28X28_x757 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x757),
 .score_0 (score_0_x757),
 .score_1 (score_1_x757),
 .score_2 (score_2_x757),
 .score_3 (score_3_x757),
 .score_4 (score_4_x757),
 .score_5 (score_5_x757),
 .score_6 (score_6_x757),
 .score_7 (score_7_x757),
 .score_8 (score_8_x757),
 .score_9 (score_9_x757)
);
 
myram_28X28 #(
.ID(758),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x758),
.W_1(W_1_x758),
.W_2(W_2_x758),
.W_3(W_3_x758),
.W_4(W_4_x758),
.W_5(W_5_x758),
.W_6(W_6_x758),
.W_7(W_7_x758),
.W_8(W_8_x758),
.W_9(W_9_x758)
) u_28X28_x758 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x758),
 .score_0 (score_0_x758),
 .score_1 (score_1_x758),
 .score_2 (score_2_x758),
 .score_3 (score_3_x758),
 .score_4 (score_4_x758),
 .score_5 (score_5_x758),
 .score_6 (score_6_x758),
 .score_7 (score_7_x758),
 .score_8 (score_8_x758),
 .score_9 (score_9_x758)
);
 
myram_28X28 #(
.ID(759),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x759),
.W_1(W_1_x759),
.W_2(W_2_x759),
.W_3(W_3_x759),
.W_4(W_4_x759),
.W_5(W_5_x759),
.W_6(W_6_x759),
.W_7(W_7_x759),
.W_8(W_8_x759),
.W_9(W_9_x759)
) u_28X28_x759 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x759),
 .score_0 (score_0_x759),
 .score_1 (score_1_x759),
 .score_2 (score_2_x759),
 .score_3 (score_3_x759),
 .score_4 (score_4_x759),
 .score_5 (score_5_x759),
 .score_6 (score_6_x759),
 .score_7 (score_7_x759),
 .score_8 (score_8_x759),
 .score_9 (score_9_x759)
);
 
myram_28X28 #(
.ID(760),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x760),
.W_1(W_1_x760),
.W_2(W_2_x760),
.W_3(W_3_x760),
.W_4(W_4_x760),
.W_5(W_5_x760),
.W_6(W_6_x760),
.W_7(W_7_x760),
.W_8(W_8_x760),
.W_9(W_9_x760)
) u_28X28_x760 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x760),
 .score_0 (score_0_x760),
 .score_1 (score_1_x760),
 .score_2 (score_2_x760),
 .score_3 (score_3_x760),
 .score_4 (score_4_x760),
 .score_5 (score_5_x760),
 .score_6 (score_6_x760),
 .score_7 (score_7_x760),
 .score_8 (score_8_x760),
 .score_9 (score_9_x760)
);
 
myram_28X28 #(
.ID(761),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x761),
.W_1(W_1_x761),
.W_2(W_2_x761),
.W_3(W_3_x761),
.W_4(W_4_x761),
.W_5(W_5_x761),
.W_6(W_6_x761),
.W_7(W_7_x761),
.W_8(W_8_x761),
.W_9(W_9_x761)
) u_28X28_x761 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x761),
 .score_0 (score_0_x761),
 .score_1 (score_1_x761),
 .score_2 (score_2_x761),
 .score_3 (score_3_x761),
 .score_4 (score_4_x761),
 .score_5 (score_5_x761),
 .score_6 (score_6_x761),
 .score_7 (score_7_x761),
 .score_8 (score_8_x761),
 .score_9 (score_9_x761)
);
 
myram_28X28 #(
.ID(762),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x762),
.W_1(W_1_x762),
.W_2(W_2_x762),
.W_3(W_3_x762),
.W_4(W_4_x762),
.W_5(W_5_x762),
.W_6(W_6_x762),
.W_7(W_7_x762),
.W_8(W_8_x762),
.W_9(W_9_x762)
) u_28X28_x762 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x762),
 .score_0 (score_0_x762),
 .score_1 (score_1_x762),
 .score_2 (score_2_x762),
 .score_3 (score_3_x762),
 .score_4 (score_4_x762),
 .score_5 (score_5_x762),
 .score_6 (score_6_x762),
 .score_7 (score_7_x762),
 .score_8 (score_8_x762),
 .score_9 (score_9_x762)
);
 
myram_28X28 #(
.ID(763),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x763),
.W_1(W_1_x763),
.W_2(W_2_x763),
.W_3(W_3_x763),
.W_4(W_4_x763),
.W_5(W_5_x763),
.W_6(W_6_x763),
.W_7(W_7_x763),
.W_8(W_8_x763),
.W_9(W_9_x763)
) u_28X28_x763 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x763),
 .score_0 (score_0_x763),
 .score_1 (score_1_x763),
 .score_2 (score_2_x763),
 .score_3 (score_3_x763),
 .score_4 (score_4_x763),
 .score_5 (score_5_x763),
 .score_6 (score_6_x763),
 .score_7 (score_7_x763),
 .score_8 (score_8_x763),
 .score_9 (score_9_x763)
);
 
myram_28X28 #(
.ID(764),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x764),
.W_1(W_1_x764),
.W_2(W_2_x764),
.W_3(W_3_x764),
.W_4(W_4_x764),
.W_5(W_5_x764),
.W_6(W_6_x764),
.W_7(W_7_x764),
.W_8(W_8_x764),
.W_9(W_9_x764)
) u_28X28_x764 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x764),
 .score_0 (score_0_x764),
 .score_1 (score_1_x764),
 .score_2 (score_2_x764),
 .score_3 (score_3_x764),
 .score_4 (score_4_x764),
 .score_5 (score_5_x764),
 .score_6 (score_6_x764),
 .score_7 (score_7_x764),
 .score_8 (score_8_x764),
 .score_9 (score_9_x764)
);
 
myram_28X28 #(
.ID(765),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x765),
.W_1(W_1_x765),
.W_2(W_2_x765),
.W_3(W_3_x765),
.W_4(W_4_x765),
.W_5(W_5_x765),
.W_6(W_6_x765),
.W_7(W_7_x765),
.W_8(W_8_x765),
.W_9(W_9_x765)
) u_28X28_x765 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x765),
 .score_0 (score_0_x765),
 .score_1 (score_1_x765),
 .score_2 (score_2_x765),
 .score_3 (score_3_x765),
 .score_4 (score_4_x765),
 .score_5 (score_5_x765),
 .score_6 (score_6_x765),
 .score_7 (score_7_x765),
 .score_8 (score_8_x765),
 .score_9 (score_9_x765)
);
 
myram_28X28 #(
.ID(766),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x766),
.W_1(W_1_x766),
.W_2(W_2_x766),
.W_3(W_3_x766),
.W_4(W_4_x766),
.W_5(W_5_x766),
.W_6(W_6_x766),
.W_7(W_7_x766),
.W_8(W_8_x766),
.W_9(W_9_x766)
) u_28X28_x766 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x766),
 .score_0 (score_0_x766),
 .score_1 (score_1_x766),
 .score_2 (score_2_x766),
 .score_3 (score_3_x766),
 .score_4 (score_4_x766),
 .score_5 (score_5_x766),
 .score_6 (score_6_x766),
 .score_7 (score_7_x766),
 .score_8 (score_8_x766),
 .score_9 (score_9_x766)
);
 
myram_28X28 #(
.ID(767),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x767),
.W_1(W_1_x767),
.W_2(W_2_x767),
.W_3(W_3_x767),
.W_4(W_4_x767),
.W_5(W_5_x767),
.W_6(W_6_x767),
.W_7(W_7_x767),
.W_8(W_8_x767),
.W_9(W_9_x767)
) u_28X28_x767 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x767),
 .score_0 (score_0_x767),
 .score_1 (score_1_x767),
 .score_2 (score_2_x767),
 .score_3 (score_3_x767),
 .score_4 (score_4_x767),
 .score_5 (score_5_x767),
 .score_6 (score_6_x767),
 .score_7 (score_7_x767),
 .score_8 (score_8_x767),
 .score_9 (score_9_x767)
);
 
myram_28X28 #(
.ID(768),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x768),
.W_1(W_1_x768),
.W_2(W_2_x768),
.W_3(W_3_x768),
.W_4(W_4_x768),
.W_5(W_5_x768),
.W_6(W_6_x768),
.W_7(W_7_x768),
.W_8(W_8_x768),
.W_9(W_9_x768)
) u_28X28_x768 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x768),
 .score_0 (score_0_x768),
 .score_1 (score_1_x768),
 .score_2 (score_2_x768),
 .score_3 (score_3_x768),
 .score_4 (score_4_x768),
 .score_5 (score_5_x768),
 .score_6 (score_6_x768),
 .score_7 (score_7_x768),
 .score_8 (score_8_x768),
 .score_9 (score_9_x768)
);
 
myram_28X28 #(
.ID(769),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x769),
.W_1(W_1_x769),
.W_2(W_2_x769),
.W_3(W_3_x769),
.W_4(W_4_x769),
.W_5(W_5_x769),
.W_6(W_6_x769),
.W_7(W_7_x769),
.W_8(W_8_x769),
.W_9(W_9_x769)
) u_28X28_x769 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x769),
 .score_0 (score_0_x769),
 .score_1 (score_1_x769),
 .score_2 (score_2_x769),
 .score_3 (score_3_x769),
 .score_4 (score_4_x769),
 .score_5 (score_5_x769),
 .score_6 (score_6_x769),
 .score_7 (score_7_x769),
 .score_8 (score_8_x769),
 .score_9 (score_9_x769)
);
 
myram_28X28 #(
.ID(770),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x770),
.W_1(W_1_x770),
.W_2(W_2_x770),
.W_3(W_3_x770),
.W_4(W_4_x770),
.W_5(W_5_x770),
.W_6(W_6_x770),
.W_7(W_7_x770),
.W_8(W_8_x770),
.W_9(W_9_x770)
) u_28X28_x770 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x770),
 .score_0 (score_0_x770),
 .score_1 (score_1_x770),
 .score_2 (score_2_x770),
 .score_3 (score_3_x770),
 .score_4 (score_4_x770),
 .score_5 (score_5_x770),
 .score_6 (score_6_x770),
 .score_7 (score_7_x770),
 .score_8 (score_8_x770),
 .score_9 (score_9_x770)
);
 
myram_28X28 #(
.ID(771),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x771),
.W_1(W_1_x771),
.W_2(W_2_x771),
.W_3(W_3_x771),
.W_4(W_4_x771),
.W_5(W_5_x771),
.W_6(W_6_x771),
.W_7(W_7_x771),
.W_8(W_8_x771),
.W_9(W_9_x771)
) u_28X28_x771 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x771),
 .score_0 (score_0_x771),
 .score_1 (score_1_x771),
 .score_2 (score_2_x771),
 .score_3 (score_3_x771),
 .score_4 (score_4_x771),
 .score_5 (score_5_x771),
 .score_6 (score_6_x771),
 .score_7 (score_7_x771),
 .score_8 (score_8_x771),
 .score_9 (score_9_x771)
);
 
myram_28X28 #(
.ID(772),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x772),
.W_1(W_1_x772),
.W_2(W_2_x772),
.W_3(W_3_x772),
.W_4(W_4_x772),
.W_5(W_5_x772),
.W_6(W_6_x772),
.W_7(W_7_x772),
.W_8(W_8_x772),
.W_9(W_9_x772)
) u_28X28_x772 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x772),
 .score_0 (score_0_x772),
 .score_1 (score_1_x772),
 .score_2 (score_2_x772),
 .score_3 (score_3_x772),
 .score_4 (score_4_x772),
 .score_5 (score_5_x772),
 .score_6 (score_6_x772),
 .score_7 (score_7_x772),
 .score_8 (score_8_x772),
 .score_9 (score_9_x772)
);
 
myram_28X28 #(
.ID(773),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x773),
.W_1(W_1_x773),
.W_2(W_2_x773),
.W_3(W_3_x773),
.W_4(W_4_x773),
.W_5(W_5_x773),
.W_6(W_6_x773),
.W_7(W_7_x773),
.W_8(W_8_x773),
.W_9(W_9_x773)
) u_28X28_x773 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x773),
 .score_0 (score_0_x773),
 .score_1 (score_1_x773),
 .score_2 (score_2_x773),
 .score_3 (score_3_x773),
 .score_4 (score_4_x773),
 .score_5 (score_5_x773),
 .score_6 (score_6_x773),
 .score_7 (score_7_x773),
 .score_8 (score_8_x773),
 .score_9 (score_9_x773)
);
 
myram_28X28 #(
.ID(774),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x774),
.W_1(W_1_x774),
.W_2(W_2_x774),
.W_3(W_3_x774),
.W_4(W_4_x774),
.W_5(W_5_x774),
.W_6(W_6_x774),
.W_7(W_7_x774),
.W_8(W_8_x774),
.W_9(W_9_x774)
) u_28X28_x774 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x774),
 .score_0 (score_0_x774),
 .score_1 (score_1_x774),
 .score_2 (score_2_x774),
 .score_3 (score_3_x774),
 .score_4 (score_4_x774),
 .score_5 (score_5_x774),
 .score_6 (score_6_x774),
 .score_7 (score_7_x774),
 .score_8 (score_8_x774),
 .score_9 (score_9_x774)
);
 
myram_28X28 #(
.ID(775),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x775),
.W_1(W_1_x775),
.W_2(W_2_x775),
.W_3(W_3_x775),
.W_4(W_4_x775),
.W_5(W_5_x775),
.W_6(W_6_x775),
.W_7(W_7_x775),
.W_8(W_8_x775),
.W_9(W_9_x775)
) u_28X28_x775 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x775),
 .score_0 (score_0_x775),
 .score_1 (score_1_x775),
 .score_2 (score_2_x775),
 .score_3 (score_3_x775),
 .score_4 (score_4_x775),
 .score_5 (score_5_x775),
 .score_6 (score_6_x775),
 .score_7 (score_7_x775),
 .score_8 (score_8_x775),
 .score_9 (score_9_x775)
);
 
myram_28X28 #(
.ID(776),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x776),
.W_1(W_1_x776),
.W_2(W_2_x776),
.W_3(W_3_x776),
.W_4(W_4_x776),
.W_5(W_5_x776),
.W_6(W_6_x776),
.W_7(W_7_x776),
.W_8(W_8_x776),
.W_9(W_9_x776)
) u_28X28_x776 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x776),
 .score_0 (score_0_x776),
 .score_1 (score_1_x776),
 .score_2 (score_2_x776),
 .score_3 (score_3_x776),
 .score_4 (score_4_x776),
 .score_5 (score_5_x776),
 .score_6 (score_6_x776),
 .score_7 (score_7_x776),
 .score_8 (score_8_x776),
 .score_9 (score_9_x776)
);
 
myram_28X28 #(
.ID(777),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x777),
.W_1(W_1_x777),
.W_2(W_2_x777),
.W_3(W_3_x777),
.W_4(W_4_x777),
.W_5(W_5_x777),
.W_6(W_6_x777),
.W_7(W_7_x777),
.W_8(W_8_x777),
.W_9(W_9_x777)
) u_28X28_x777 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x777),
 .score_0 (score_0_x777),
 .score_1 (score_1_x777),
 .score_2 (score_2_x777),
 .score_3 (score_3_x777),
 .score_4 (score_4_x777),
 .score_5 (score_5_x777),
 .score_6 (score_6_x777),
 .score_7 (score_7_x777),
 .score_8 (score_8_x777),
 .score_9 (score_9_x777)
);
 
myram_28X28 #(
.ID(778),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x778),
.W_1(W_1_x778),
.W_2(W_2_x778),
.W_3(W_3_x778),
.W_4(W_4_x778),
.W_5(W_5_x778),
.W_6(W_6_x778),
.W_7(W_7_x778),
.W_8(W_8_x778),
.W_9(W_9_x778)
) u_28X28_x778 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x778),
 .score_0 (score_0_x778),
 .score_1 (score_1_x778),
 .score_2 (score_2_x778),
 .score_3 (score_3_x778),
 .score_4 (score_4_x778),
 .score_5 (score_5_x778),
 .score_6 (score_6_x778),
 .score_7 (score_7_x778),
 .score_8 (score_8_x778),
 .score_9 (score_9_x778)
);
 
myram_28X28 #(
.ID(779),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x779),
.W_1(W_1_x779),
.W_2(W_2_x779),
.W_3(W_3_x779),
.W_4(W_4_x779),
.W_5(W_5_x779),
.W_6(W_6_x779),
.W_7(W_7_x779),
.W_8(W_8_x779),
.W_9(W_9_x779)
) u_28X28_x779 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x779),
 .score_0 (score_0_x779),
 .score_1 (score_1_x779),
 .score_2 (score_2_x779),
 .score_3 (score_3_x779),
 .score_4 (score_4_x779),
 .score_5 (score_5_x779),
 .score_6 (score_6_x779),
 .score_7 (score_7_x779),
 .score_8 (score_8_x779),
 .score_9 (score_9_x779)
);
 
myram_28X28 #(
.ID(780),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x780),
.W_1(W_1_x780),
.W_2(W_2_x780),
.W_3(W_3_x780),
.W_4(W_4_x780),
.W_5(W_5_x780),
.W_6(W_6_x780),
.W_7(W_7_x780),
.W_8(W_8_x780),
.W_9(W_9_x780)
) u_28X28_x780 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x780),
 .score_0 (score_0_x780),
 .score_1 (score_1_x780),
 .score_2 (score_2_x780),
 .score_3 (score_3_x780),
 .score_4 (score_4_x780),
 .score_5 (score_5_x780),
 .score_6 (score_6_x780),
 .score_7 (score_7_x780),
 .score_8 (score_8_x780),
 .score_9 (score_9_x780)
);
 
myram_28X28 #(
.ID(781),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x781),
.W_1(W_1_x781),
.W_2(W_2_x781),
.W_3(W_3_x781),
.W_4(W_4_x781),
.W_5(W_5_x781),
.W_6(W_6_x781),
.W_7(W_7_x781),
.W_8(W_8_x781),
.W_9(W_9_x781)
) u_28X28_x781 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x781),
 .score_0 (score_0_x781),
 .score_1 (score_1_x781),
 .score_2 (score_2_x781),
 .score_3 (score_3_x781),
 .score_4 (score_4_x781),
 .score_5 (score_5_x781),
 .score_6 (score_6_x781),
 .score_7 (score_7_x781),
 .score_8 (score_8_x781),
 .score_9 (score_9_x781)
);
 
myram_28X28 #(
.ID(782),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x782),
.W_1(W_1_x782),
.W_2(W_2_x782),
.W_3(W_3_x782),
.W_4(W_4_x782),
.W_5(W_5_x782),
.W_6(W_6_x782),
.W_7(W_7_x782),
.W_8(W_8_x782),
.W_9(W_9_x782)
) u_28X28_x782 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x782),
 .score_0 (score_0_x782),
 .score_1 (score_1_x782),
 .score_2 (score_2_x782),
 .score_3 (score_3_x782),
 .score_4 (score_4_x782),
 .score_5 (score_5_x782),
 .score_6 (score_6_x782),
 .score_7 (score_7_x782),
 .score_8 (score_8_x782),
 .score_9 (score_9_x782)
);
 
myram_28X28 #(
.ID(783),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x783),
.W_1(W_1_x783),
.W_2(W_2_x783),
.W_3(W_3_x783),
.W_4(W_4_x783),
.W_5(W_5_x783),
.W_6(W_6_x783),
.W_7(W_7_x783),
.W_8(W_8_x783),
.W_9(W_9_x783)
) u_28X28_x783 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x783),
 .score_0 (score_0_x783),
 .score_1 (score_1_x783),
 .score_2 (score_2_x783),
 .score_3 (score_3_x783),
 .score_4 (score_4_x783),
 .score_5 (score_5_x783),
 .score_6 (score_6_x783),
 .score_7 (score_7_x783),
 .score_8 (score_8_x783),
 .score_9 (score_9_x783)
);
 
myram_28X28 #(
.ID(784),
.UP(UP),
.DOWN(DOWN),
.LEFT(LEFT),
.RIGHT(RIGHT),
.EACH_WIDE(EACH_WIDE),.DEBIT(DEBIT),
.W_0(W_0_x784),
.W_1(W_1_x784),
.W_2(W_2_x784),
.W_3(W_3_x784),
.W_4(W_4_x784),
.W_5(W_5_x784),
.W_6(W_6_x784),
.W_7(W_7_x784),
.W_8(W_8_x784),
.W_9(W_9_x784)
) u_28X28_x784 (
 .clk (clk),
 .xpos (xpos),
 .ypos (ypos),
 .dq_i (dq_i),
 .res_done (res_done_x784),
 .score_0 (score_0_x784),
 .score_1 (score_1_x784),
 .score_2 (score_2_x784),
 .score_3 (score_3_x784),
 .score_4 (score_4_x784),
 .score_5 (score_5_x784),
 .score_6 (score_6_x784),
 .score_7 (score_7_x784),
 .score_8 (score_8_x784),
 .score_9 (score_9_x784)
);
 



    
endmodule